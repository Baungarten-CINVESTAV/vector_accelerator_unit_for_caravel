// This is the unpowered netlist.
module ALU (Exception,
    Overflow,
    Underflow,
    ALU_Output,
    Operation,
    a_operand,
    b_operand);
 output Exception;
 output Overflow;
 output Underflow;
 output [31:0] ALU_Output;
 input [3:0] Operation;
 input [31:0] a_operand;
 input [31:0] b_operand;

 wire \AuI.AddBar_Sub ;
 wire \AuI.Exception ;
 wire \AuI._0000_ ;
 wire \AuI._0001_ ;
 wire \AuI._0002_ ;
 wire \AuI._0003_ ;
 wire \AuI._0004_ ;
 wire \AuI._0005_ ;
 wire \AuI._0006_ ;
 wire \AuI._0007_ ;
 wire \AuI._0008_ ;
 wire \AuI._0009_ ;
 wire \AuI._0010_ ;
 wire \AuI._0011_ ;
 wire \AuI._0012_ ;
 wire \AuI._0013_ ;
 wire \AuI._0014_ ;
 wire \AuI._0015_ ;
 wire \AuI._0016_ ;
 wire \AuI._0017_ ;
 wire \AuI._0018_ ;
 wire \AuI._0019_ ;
 wire \AuI._0020_ ;
 wire \AuI._0021_ ;
 wire \AuI._0022_ ;
 wire \AuI._0023_ ;
 wire \AuI._0024_ ;
 wire \AuI._0025_ ;
 wire \AuI._0026_ ;
 wire \AuI._0027_ ;
 wire \AuI._0028_ ;
 wire \AuI._0029_ ;
 wire \AuI._0030_ ;
 wire \AuI._0031_ ;
 wire \AuI._0032_ ;
 wire \AuI._0033_ ;
 wire \AuI._0034_ ;
 wire \AuI._0035_ ;
 wire \AuI._0036_ ;
 wire \AuI._0037_ ;
 wire \AuI._0038_ ;
 wire \AuI._0039_ ;
 wire \AuI._0040_ ;
 wire \AuI._0041_ ;
 wire \AuI._0042_ ;
 wire \AuI._0043_ ;
 wire \AuI._0044_ ;
 wire \AuI._0045_ ;
 wire \AuI._0046_ ;
 wire \AuI._0047_ ;
 wire \AuI._0048_ ;
 wire \AuI._0049_ ;
 wire \AuI._0050_ ;
 wire \AuI._0051_ ;
 wire \AuI._0052_ ;
 wire \AuI._0053_ ;
 wire \AuI._0054_ ;
 wire \AuI._0055_ ;
 wire \AuI._0056_ ;
 wire \AuI._0057_ ;
 wire \AuI._0058_ ;
 wire \AuI._0059_ ;
 wire \AuI._0060_ ;
 wire \AuI._0061_ ;
 wire \AuI._0062_ ;
 wire \AuI._0063_ ;
 wire \AuI._0064_ ;
 wire \AuI._0065_ ;
 wire \AuI._0066_ ;
 wire \AuI._0067_ ;
 wire \AuI._0068_ ;
 wire \AuI._0069_ ;
 wire \AuI._0070_ ;
 wire \AuI._0071_ ;
 wire \AuI._0072_ ;
 wire \AuI._0073_ ;
 wire \AuI._0074_ ;
 wire \AuI._0075_ ;
 wire \AuI._0076_ ;
 wire \AuI._0077_ ;
 wire \AuI._0078_ ;
 wire \AuI._0079_ ;
 wire \AuI._0080_ ;
 wire \AuI._0081_ ;
 wire \AuI._0082_ ;
 wire \AuI._0083_ ;
 wire \AuI._0084_ ;
 wire \AuI._0085_ ;
 wire \AuI._0086_ ;
 wire \AuI._0087_ ;
 wire \AuI._0088_ ;
 wire \AuI._0089_ ;
 wire \AuI._0090_ ;
 wire \AuI._0091_ ;
 wire \AuI._0092_ ;
 wire \AuI._0093_ ;
 wire \AuI._0094_ ;
 wire \AuI._0095_ ;
 wire \AuI._0096_ ;
 wire \AuI._0097_ ;
 wire \AuI._0098_ ;
 wire \AuI._0099_ ;
 wire \AuI._0100_ ;
 wire \AuI._0101_ ;
 wire \AuI._0102_ ;
 wire \AuI._0103_ ;
 wire \AuI._0104_ ;
 wire \AuI._0105_ ;
 wire \AuI._0106_ ;
 wire \AuI._0107_ ;
 wire \AuI._0108_ ;
 wire \AuI._0109_ ;
 wire \AuI._0110_ ;
 wire \AuI._0111_ ;
 wire \AuI._0112_ ;
 wire \AuI._0113_ ;
 wire \AuI._0114_ ;
 wire \AuI._0115_ ;
 wire \AuI._0116_ ;
 wire \AuI._0117_ ;
 wire \AuI._0118_ ;
 wire \AuI._0119_ ;
 wire \AuI._0120_ ;
 wire \AuI._0121_ ;
 wire \AuI._0122_ ;
 wire \AuI._0123_ ;
 wire \AuI._0124_ ;
 wire \AuI._0125_ ;
 wire \AuI._0126_ ;
 wire \AuI._0127_ ;
 wire \AuI._0128_ ;
 wire \AuI._0129_ ;
 wire \AuI._0130_ ;
 wire \AuI._0131_ ;
 wire \AuI._0132_ ;
 wire \AuI._0133_ ;
 wire \AuI._0134_ ;
 wire \AuI._0135_ ;
 wire \AuI._0136_ ;
 wire \AuI._0137_ ;
 wire \AuI._0138_ ;
 wire \AuI._0139_ ;
 wire \AuI._0140_ ;
 wire \AuI._0141_ ;
 wire \AuI._0142_ ;
 wire \AuI._0143_ ;
 wire \AuI._0144_ ;
 wire \AuI._0145_ ;
 wire \AuI._0146_ ;
 wire \AuI._0147_ ;
 wire \AuI._0148_ ;
 wire \AuI._0149_ ;
 wire \AuI._0150_ ;
 wire \AuI._0151_ ;
 wire \AuI._0152_ ;
 wire \AuI._0153_ ;
 wire \AuI._0154_ ;
 wire \AuI._0155_ ;
 wire \AuI._0156_ ;
 wire \AuI._0157_ ;
 wire \AuI._0158_ ;
 wire \AuI._0159_ ;
 wire \AuI._0160_ ;
 wire \AuI._0161_ ;
 wire \AuI._0162_ ;
 wire \AuI._0163_ ;
 wire \AuI._0164_ ;
 wire \AuI._0165_ ;
 wire \AuI._0166_ ;
 wire \AuI._0167_ ;
 wire \AuI._0168_ ;
 wire \AuI._0169_ ;
 wire \AuI._0170_ ;
 wire \AuI._0171_ ;
 wire \AuI._0172_ ;
 wire \AuI._0173_ ;
 wire \AuI._0174_ ;
 wire \AuI._0175_ ;
 wire \AuI._0176_ ;
 wire \AuI._0177_ ;
 wire \AuI._0178_ ;
 wire \AuI._0179_ ;
 wire \AuI._0180_ ;
 wire \AuI._0181_ ;
 wire \AuI._0182_ ;
 wire \AuI._0183_ ;
 wire \AuI._0184_ ;
 wire \AuI._0185_ ;
 wire \AuI._0186_ ;
 wire \AuI._0187_ ;
 wire \AuI._0188_ ;
 wire \AuI._0189_ ;
 wire \AuI._0190_ ;
 wire \AuI._0191_ ;
 wire \AuI._0192_ ;
 wire \AuI._0193_ ;
 wire \AuI._0194_ ;
 wire \AuI._0195_ ;
 wire \AuI._0196_ ;
 wire \AuI._0197_ ;
 wire \AuI._0198_ ;
 wire \AuI._0199_ ;
 wire \AuI._0200_ ;
 wire \AuI._0201_ ;
 wire \AuI._0202_ ;
 wire \AuI._0203_ ;
 wire \AuI._0204_ ;
 wire \AuI._0205_ ;
 wire \AuI._0206_ ;
 wire \AuI._0207_ ;
 wire \AuI._0208_ ;
 wire \AuI._0209_ ;
 wire \AuI._0210_ ;
 wire \AuI._0211_ ;
 wire \AuI._0212_ ;
 wire \AuI._0213_ ;
 wire \AuI._0214_ ;
 wire \AuI._0215_ ;
 wire \AuI._0216_ ;
 wire \AuI._0217_ ;
 wire \AuI._0218_ ;
 wire \AuI._0219_ ;
 wire \AuI._0220_ ;
 wire \AuI._0221_ ;
 wire \AuI._0222_ ;
 wire \AuI._0223_ ;
 wire \AuI._0224_ ;
 wire \AuI._0225_ ;
 wire \AuI._0226_ ;
 wire \AuI._0227_ ;
 wire \AuI._0228_ ;
 wire \AuI._0229_ ;
 wire \AuI._0230_ ;
 wire \AuI._0231_ ;
 wire \AuI._0232_ ;
 wire \AuI._0233_ ;
 wire \AuI._0234_ ;
 wire \AuI._0235_ ;
 wire \AuI._0236_ ;
 wire \AuI._0237_ ;
 wire \AuI._0238_ ;
 wire \AuI._0239_ ;
 wire \AuI._0240_ ;
 wire \AuI._0241_ ;
 wire \AuI._0242_ ;
 wire \AuI._0243_ ;
 wire \AuI._0244_ ;
 wire \AuI._0245_ ;
 wire \AuI._0246_ ;
 wire \AuI._0247_ ;
 wire \AuI._0248_ ;
 wire \AuI._0249_ ;
 wire \AuI._0250_ ;
 wire \AuI._0251_ ;
 wire \AuI._0252_ ;
 wire \AuI._0253_ ;
 wire \AuI._0254_ ;
 wire \AuI._0255_ ;
 wire \AuI._0256_ ;
 wire \AuI._0257_ ;
 wire \AuI._0258_ ;
 wire \AuI._0259_ ;
 wire \AuI._0260_ ;
 wire \AuI._0261_ ;
 wire \AuI._0262_ ;
 wire \AuI._0263_ ;
 wire \AuI._0264_ ;
 wire \AuI._0265_ ;
 wire \AuI._0266_ ;
 wire \AuI._0267_ ;
 wire \AuI._0268_ ;
 wire \AuI._0269_ ;
 wire \AuI._0270_ ;
 wire \AuI._0271_ ;
 wire \AuI._0272_ ;
 wire \AuI._0273_ ;
 wire \AuI._0274_ ;
 wire \AuI._0275_ ;
 wire \AuI._0276_ ;
 wire \AuI._0277_ ;
 wire \AuI._0278_ ;
 wire \AuI._0279_ ;
 wire \AuI._0280_ ;
 wire \AuI._0281_ ;
 wire \AuI._0282_ ;
 wire \AuI._0283_ ;
 wire \AuI._0284_ ;
 wire \AuI._0285_ ;
 wire \AuI._0286_ ;
 wire \AuI._0287_ ;
 wire \AuI._0288_ ;
 wire \AuI._0289_ ;
 wire \AuI._0290_ ;
 wire \AuI._0291_ ;
 wire \AuI._0292_ ;
 wire \AuI._0293_ ;
 wire \AuI._0294_ ;
 wire \AuI._0295_ ;
 wire \AuI._0296_ ;
 wire \AuI._0297_ ;
 wire \AuI._0298_ ;
 wire \AuI._0299_ ;
 wire \AuI._0300_ ;
 wire \AuI._0301_ ;
 wire \AuI._0302_ ;
 wire \AuI._0303_ ;
 wire \AuI._0304_ ;
 wire \AuI._0305_ ;
 wire \AuI._0306_ ;
 wire \AuI._0307_ ;
 wire \AuI._0308_ ;
 wire \AuI._0309_ ;
 wire \AuI._0310_ ;
 wire \AuI._0311_ ;
 wire \AuI._0312_ ;
 wire \AuI._0313_ ;
 wire \AuI._0314_ ;
 wire \AuI._0315_ ;
 wire \AuI._0316_ ;
 wire \AuI._0317_ ;
 wire \AuI._0318_ ;
 wire \AuI._0319_ ;
 wire \AuI._0320_ ;
 wire \AuI._0321_ ;
 wire \AuI._0322_ ;
 wire \AuI._0323_ ;
 wire \AuI._0324_ ;
 wire \AuI._0325_ ;
 wire \AuI._0326_ ;
 wire \AuI._0327_ ;
 wire \AuI._0328_ ;
 wire \AuI._0329_ ;
 wire \AuI._0330_ ;
 wire \AuI._0331_ ;
 wire \AuI._0332_ ;
 wire \AuI._0333_ ;
 wire \AuI._0334_ ;
 wire \AuI._0335_ ;
 wire \AuI._0336_ ;
 wire \AuI._0337_ ;
 wire \AuI._0338_ ;
 wire \AuI._0339_ ;
 wire \AuI._0340_ ;
 wire \AuI._0341_ ;
 wire \AuI._0342_ ;
 wire \AuI._0343_ ;
 wire \AuI._0344_ ;
 wire \AuI._0345_ ;
 wire \AuI._0346_ ;
 wire \AuI._0347_ ;
 wire \AuI._0348_ ;
 wire \AuI._0349_ ;
 wire \AuI._0350_ ;
 wire \AuI._0351_ ;
 wire \AuI._0352_ ;
 wire \AuI._0353_ ;
 wire \AuI._0354_ ;
 wire \AuI._0355_ ;
 wire \AuI._0356_ ;
 wire \AuI._0357_ ;
 wire \AuI._0358_ ;
 wire \AuI._0359_ ;
 wire \AuI._0360_ ;
 wire \AuI._0361_ ;
 wire \AuI._0362_ ;
 wire \AuI._0363_ ;
 wire \AuI._0364_ ;
 wire \AuI._0365_ ;
 wire \AuI._0366_ ;
 wire \AuI._0367_ ;
 wire \AuI._0368_ ;
 wire \AuI._0369_ ;
 wire \AuI._0370_ ;
 wire \AuI._0371_ ;
 wire \AuI._0372_ ;
 wire \AuI._0373_ ;
 wire \AuI._0374_ ;
 wire \AuI._0375_ ;
 wire \AuI._0376_ ;
 wire \AuI._0377_ ;
 wire \AuI._0378_ ;
 wire \AuI._0379_ ;
 wire \AuI._0380_ ;
 wire \AuI._0381_ ;
 wire \AuI._0382_ ;
 wire \AuI._0383_ ;
 wire \AuI._0384_ ;
 wire \AuI._0385_ ;
 wire \AuI._0386_ ;
 wire \AuI._0387_ ;
 wire \AuI._0388_ ;
 wire \AuI._0389_ ;
 wire \AuI._0390_ ;
 wire \AuI._0391_ ;
 wire \AuI._0392_ ;
 wire \AuI._0393_ ;
 wire \AuI._0394_ ;
 wire \AuI._0395_ ;
 wire \AuI._0396_ ;
 wire \AuI._0397_ ;
 wire \AuI._0398_ ;
 wire \AuI._0399_ ;
 wire \AuI._0400_ ;
 wire \AuI._0401_ ;
 wire \AuI._0402_ ;
 wire \AuI._0403_ ;
 wire \AuI._0404_ ;
 wire \AuI._0405_ ;
 wire \AuI._0406_ ;
 wire \AuI._0407_ ;
 wire \AuI._0408_ ;
 wire \AuI._0409_ ;
 wire \AuI._0410_ ;
 wire \AuI._0411_ ;
 wire \AuI._0412_ ;
 wire \AuI._0413_ ;
 wire \AuI._0414_ ;
 wire \AuI._0415_ ;
 wire \AuI._0416_ ;
 wire \AuI._0417_ ;
 wire \AuI._0418_ ;
 wire \AuI._0419_ ;
 wire \AuI._0420_ ;
 wire \AuI._0421_ ;
 wire \AuI._0422_ ;
 wire \AuI._0423_ ;
 wire \AuI._0424_ ;
 wire \AuI._0425_ ;
 wire \AuI._0426_ ;
 wire \AuI._0427_ ;
 wire \AuI._0428_ ;
 wire \AuI._0429_ ;
 wire \AuI._0430_ ;
 wire \AuI._0431_ ;
 wire \AuI._0432_ ;
 wire \AuI._0433_ ;
 wire \AuI._0434_ ;
 wire \AuI._0435_ ;
 wire \AuI._0436_ ;
 wire \AuI._0437_ ;
 wire \AuI._0438_ ;
 wire \AuI._0439_ ;
 wire \AuI._0440_ ;
 wire \AuI._0441_ ;
 wire \AuI._0442_ ;
 wire \AuI._0443_ ;
 wire \AuI._0444_ ;
 wire \AuI._0445_ ;
 wire \AuI._0446_ ;
 wire \AuI._0447_ ;
 wire \AuI._0448_ ;
 wire \AuI._0449_ ;
 wire \AuI._0450_ ;
 wire \AuI._0451_ ;
 wire \AuI._0452_ ;
 wire \AuI._0453_ ;
 wire \AuI._0454_ ;
 wire \AuI._0455_ ;
 wire \AuI._0456_ ;
 wire \AuI._0457_ ;
 wire \AuI._0458_ ;
 wire \AuI._0459_ ;
 wire \AuI._0460_ ;
 wire \AuI._0461_ ;
 wire \AuI._0462_ ;
 wire \AuI._0463_ ;
 wire \AuI._0464_ ;
 wire \AuI._0465_ ;
 wire \AuI._0466_ ;
 wire \AuI._0467_ ;
 wire \AuI._0468_ ;
 wire \AuI._0469_ ;
 wire \AuI._0470_ ;
 wire \AuI._0471_ ;
 wire \AuI._0472_ ;
 wire \AuI._0473_ ;
 wire \AuI._0474_ ;
 wire \AuI._0475_ ;
 wire \AuI._0476_ ;
 wire \AuI._0477_ ;
 wire \AuI._0478_ ;
 wire \AuI._0479_ ;
 wire \AuI._0480_ ;
 wire \AuI._0481_ ;
 wire \AuI._0482_ ;
 wire \AuI._0483_ ;
 wire \AuI._0484_ ;
 wire \AuI._0485_ ;
 wire \AuI._0486_ ;
 wire \AuI._0487_ ;
 wire \AuI._0488_ ;
 wire \AuI._0489_ ;
 wire \AuI._0490_ ;
 wire \AuI._0491_ ;
 wire \AuI._0492_ ;
 wire \AuI._0493_ ;
 wire \AuI._0494_ ;
 wire \AuI._0495_ ;
 wire \AuI._0496_ ;
 wire \AuI._0497_ ;
 wire \AuI._0498_ ;
 wire \AuI._0499_ ;
 wire \AuI._0500_ ;
 wire \AuI._0501_ ;
 wire \AuI._0502_ ;
 wire \AuI._0503_ ;
 wire \AuI._0504_ ;
 wire \AuI._0505_ ;
 wire \AuI._0506_ ;
 wire \AuI._0507_ ;
 wire \AuI._0508_ ;
 wire \AuI._0509_ ;
 wire \AuI._0510_ ;
 wire \AuI._0511_ ;
 wire \AuI._0512_ ;
 wire \AuI._0513_ ;
 wire \AuI._0514_ ;
 wire \AuI._0515_ ;
 wire \AuI._0516_ ;
 wire \AuI._0517_ ;
 wire \AuI._0518_ ;
 wire \AuI._0519_ ;
 wire \AuI._0520_ ;
 wire \AuI._0521_ ;
 wire \AuI._0522_ ;
 wire \AuI._0523_ ;
 wire \AuI._0524_ ;
 wire \AuI._0525_ ;
 wire \AuI._0526_ ;
 wire \AuI._0527_ ;
 wire \AuI._0528_ ;
 wire \AuI._0529_ ;
 wire \AuI._0530_ ;
 wire \AuI._0531_ ;
 wire \AuI._0532_ ;
 wire \AuI._0533_ ;
 wire \AuI._0534_ ;
 wire \AuI._0535_ ;
 wire \AuI._0536_ ;
 wire \AuI._0537_ ;
 wire \AuI._0538_ ;
 wire \AuI._0539_ ;
 wire \AuI._0540_ ;
 wire \AuI._0541_ ;
 wire \AuI._0542_ ;
 wire \AuI._0543_ ;
 wire \AuI._0544_ ;
 wire \AuI._0545_ ;
 wire \AuI._0546_ ;
 wire \AuI._0547_ ;
 wire \AuI._0548_ ;
 wire \AuI._0549_ ;
 wire \AuI._0550_ ;
 wire \AuI._0551_ ;
 wire \AuI._0552_ ;
 wire \AuI._0553_ ;
 wire \AuI._0554_ ;
 wire \AuI._0555_ ;
 wire \AuI._0556_ ;
 wire \AuI._0557_ ;
 wire \AuI._0558_ ;
 wire \AuI._0559_ ;
 wire \AuI._0560_ ;
 wire \AuI._0561_ ;
 wire \AuI._0562_ ;
 wire \AuI._0563_ ;
 wire \AuI._0564_ ;
 wire \AuI._0565_ ;
 wire \AuI._0566_ ;
 wire \AuI._0567_ ;
 wire \AuI._0568_ ;
 wire \AuI._0569_ ;
 wire \AuI._0570_ ;
 wire \AuI._0571_ ;
 wire \AuI._0572_ ;
 wire \AuI._0573_ ;
 wire \AuI._0574_ ;
 wire \AuI._0575_ ;
 wire \AuI._0576_ ;
 wire \AuI._0577_ ;
 wire \AuI._0578_ ;
 wire \AuI._0579_ ;
 wire \AuI._0580_ ;
 wire \AuI._0581_ ;
 wire \AuI._0582_ ;
 wire \AuI._0583_ ;
 wire \AuI._0584_ ;
 wire \AuI._0585_ ;
 wire \AuI._0586_ ;
 wire \AuI._0587_ ;
 wire \AuI._0588_ ;
 wire \AuI._0589_ ;
 wire \AuI._0590_ ;
 wire \AuI._0591_ ;
 wire \AuI._0592_ ;
 wire \AuI._0593_ ;
 wire \AuI._0594_ ;
 wire \AuI._0595_ ;
 wire \AuI._0596_ ;
 wire \AuI._0597_ ;
 wire \AuI._0598_ ;
 wire \AuI._0599_ ;
 wire \AuI._0600_ ;
 wire \AuI._0601_ ;
 wire \AuI._0602_ ;
 wire \AuI._0603_ ;
 wire \AuI._0604_ ;
 wire \AuI._0605_ ;
 wire \AuI._0606_ ;
 wire \AuI._0607_ ;
 wire \AuI._0608_ ;
 wire \AuI._0609_ ;
 wire \AuI._0610_ ;
 wire \AuI._0611_ ;
 wire \AuI._0612_ ;
 wire \AuI._0613_ ;
 wire \AuI._0614_ ;
 wire \AuI._0615_ ;
 wire \AuI._0616_ ;
 wire \AuI._0617_ ;
 wire \AuI._0618_ ;
 wire \AuI._0619_ ;
 wire \AuI._0620_ ;
 wire \AuI._0621_ ;
 wire \AuI._0622_ ;
 wire \AuI._0623_ ;
 wire \AuI._0624_ ;
 wire \AuI._0625_ ;
 wire \AuI._0626_ ;
 wire \AuI._0627_ ;
 wire \AuI._0628_ ;
 wire \AuI._0629_ ;
 wire \AuI._0630_ ;
 wire \AuI._0631_ ;
 wire \AuI._0632_ ;
 wire \AuI._0633_ ;
 wire \AuI._0634_ ;
 wire \AuI._0635_ ;
 wire \AuI._0636_ ;
 wire \AuI._0637_ ;
 wire \AuI._0638_ ;
 wire \AuI._0639_ ;
 wire \AuI._0640_ ;
 wire \AuI._0641_ ;
 wire \AuI._0642_ ;
 wire \AuI._0643_ ;
 wire \AuI._0644_ ;
 wire \AuI._0645_ ;
 wire \AuI._0646_ ;
 wire \AuI._0647_ ;
 wire \AuI._0648_ ;
 wire \AuI._0649_ ;
 wire \AuI._0650_ ;
 wire \AuI._0651_ ;
 wire \AuI._0652_ ;
 wire \AuI._0653_ ;
 wire \AuI._0654_ ;
 wire \AuI._0655_ ;
 wire \AuI._0656_ ;
 wire \AuI._0657_ ;
 wire \AuI._0658_ ;
 wire \AuI._0659_ ;
 wire \AuI._0660_ ;
 wire \AuI._0661_ ;
 wire \AuI._0662_ ;
 wire \AuI._0663_ ;
 wire \AuI._0664_ ;
 wire \AuI._0665_ ;
 wire \AuI._0666_ ;
 wire \AuI._0667_ ;
 wire \AuI._0668_ ;
 wire \AuI._0669_ ;
 wire \AuI._0670_ ;
 wire \AuI._0671_ ;
 wire \AuI._0672_ ;
 wire \AuI._0673_ ;
 wire \AuI._0674_ ;
 wire \AuI._0675_ ;
 wire \AuI._0676_ ;
 wire \AuI._0677_ ;
 wire \AuI._0678_ ;
 wire \AuI._0679_ ;
 wire \AuI._0680_ ;
 wire \AuI._0681_ ;
 wire \AuI._0682_ ;
 wire \AuI._0683_ ;
 wire \AuI._0684_ ;
 wire \AuI._0685_ ;
 wire \AuI._0686_ ;
 wire \AuI._0687_ ;
 wire \AuI._0688_ ;
 wire \AuI._0689_ ;
 wire \AuI._0690_ ;
 wire \AuI._0691_ ;
 wire \AuI._0692_ ;
 wire \AuI._0693_ ;
 wire \AuI._0694_ ;
 wire \AuI._0695_ ;
 wire \AuI._0696_ ;
 wire \AuI._0697_ ;
 wire \AuI._0698_ ;
 wire \AuI._0699_ ;
 wire \AuI._0700_ ;
 wire \AuI._0701_ ;
 wire \AuI._0702_ ;
 wire \AuI._0703_ ;
 wire \AuI._0704_ ;
 wire \AuI._0705_ ;
 wire \AuI._0706_ ;
 wire \AuI._0707_ ;
 wire \AuI._0708_ ;
 wire \AuI._0709_ ;
 wire \AuI._0710_ ;
 wire \AuI._0711_ ;
 wire \AuI._0712_ ;
 wire \AuI._0713_ ;
 wire \AuI._0714_ ;
 wire \AuI._0715_ ;
 wire \AuI._0716_ ;
 wire \AuI._0717_ ;
 wire \AuI._0718_ ;
 wire \AuI._0719_ ;
 wire \AuI._0720_ ;
 wire \AuI._0721_ ;
 wire \AuI._0722_ ;
 wire \AuI._0723_ ;
 wire \AuI._0724_ ;
 wire \AuI._0725_ ;
 wire \AuI._0726_ ;
 wire \AuI._0727_ ;
 wire \AuI._0728_ ;
 wire \AuI._0729_ ;
 wire \AuI._0730_ ;
 wire \AuI._0731_ ;
 wire \AuI._0732_ ;
 wire \AuI._0733_ ;
 wire \AuI._0734_ ;
 wire \AuI._0735_ ;
 wire \AuI._0736_ ;
 wire \AuI._0737_ ;
 wire \AuI._0738_ ;
 wire \AuI._0739_ ;
 wire \AuI._0740_ ;
 wire \AuI._0741_ ;
 wire \AuI._0742_ ;
 wire \AuI._0743_ ;
 wire \AuI._0744_ ;
 wire \AuI._0745_ ;
 wire \AuI._0746_ ;
 wire \AuI._0747_ ;
 wire \AuI._0748_ ;
 wire \AuI._0749_ ;
 wire \AuI._0750_ ;
 wire \AuI._0751_ ;
 wire \AuI._0752_ ;
 wire \AuI._0753_ ;
 wire \AuI._0754_ ;
 wire \AuI._0755_ ;
 wire \AuI._0756_ ;
 wire \AuI._0757_ ;
 wire \AuI._0758_ ;
 wire \AuI._0759_ ;
 wire \AuI._0760_ ;
 wire \AuI._0761_ ;
 wire \AuI._0762_ ;
 wire \AuI._0763_ ;
 wire \AuI._0764_ ;
 wire \AuI._0765_ ;
 wire \AuI._0766_ ;
 wire \AuI._0767_ ;
 wire \AuI._0768_ ;
 wire \AuI._0769_ ;
 wire \AuI._0770_ ;
 wire \AuI._0771_ ;
 wire \AuI._0772_ ;
 wire \AuI._0773_ ;
 wire \AuI._0774_ ;
 wire \AuI._0775_ ;
 wire \AuI._0776_ ;
 wire \AuI._0777_ ;
 wire \AuI._0778_ ;
 wire \AuI._0779_ ;
 wire \AuI._0780_ ;
 wire \AuI._0781_ ;
 wire \AuI._0782_ ;
 wire \AuI._0783_ ;
 wire \AuI._0784_ ;
 wire \AuI._0785_ ;
 wire \AuI._0786_ ;
 wire \AuI._0787_ ;
 wire \AuI._0788_ ;
 wire \AuI._0789_ ;
 wire \AuI._0790_ ;
 wire \AuI._0791_ ;
 wire \AuI._0792_ ;
 wire \AuI._0793_ ;
 wire \AuI._0794_ ;
 wire \AuI._0795_ ;
 wire \AuI._0796_ ;
 wire \AuI._0797_ ;
 wire \AuI._0798_ ;
 wire \AuI._0799_ ;
 wire \AuI._0800_ ;
 wire \AuI._0801_ ;
 wire \AuI._0802_ ;
 wire \AuI._0803_ ;
 wire \AuI._0804_ ;
 wire \AuI.exp_a ;
 wire \AuI.exponent_sub[0] ;
 wire \AuI.exponent_sub[1] ;
 wire \AuI.exponent_sub[2] ;
 wire \AuI.exponent_sub[3] ;
 wire \AuI.exponent_sub[4] ;
 wire \AuI.exponent_sub[5] ;
 wire \AuI.exponent_sub[6] ;
 wire \AuI.exponent_sub[7] ;
 wire \AuI.operand_a[24] ;
 wire \AuI.operand_a[25] ;
 wire \AuI.operand_a[26] ;
 wire \AuI.operand_a[27] ;
 wire \AuI.operand_a[28] ;
 wire \AuI.operand_a[29] ;
 wire \AuI.operand_a[30] ;
 wire \AuI.pe.Significand[0] ;
 wire \AuI.pe.Significand[10] ;
 wire \AuI.pe.Significand[11] ;
 wire \AuI.pe.Significand[12] ;
 wire \AuI.pe.Significand[13] ;
 wire \AuI.pe.Significand[14] ;
 wire \AuI.pe.Significand[15] ;
 wire \AuI.pe.Significand[16] ;
 wire \AuI.pe.Significand[17] ;
 wire \AuI.pe.Significand[18] ;
 wire \AuI.pe.Significand[19] ;
 wire \AuI.pe.Significand[1] ;
 wire \AuI.pe.Significand[20] ;
 wire \AuI.pe.Significand[21] ;
 wire \AuI.pe.Significand[22] ;
 wire \AuI.pe.Significand[2] ;
 wire \AuI.pe.Significand[3] ;
 wire \AuI.pe.Significand[4] ;
 wire \AuI.pe.Significand[5] ;
 wire \AuI.pe.Significand[6] ;
 wire \AuI.pe.Significand[7] ;
 wire \AuI.pe.Significand[8] ;
 wire \AuI.pe.Significand[9] ;
 wire \AuI.pe._000_ ;
 wire \AuI.pe._001_ ;
 wire \AuI.pe._002_ ;
 wire \AuI.pe._003_ ;
 wire \AuI.pe._004_ ;
 wire \AuI.pe._005_ ;
 wire \AuI.pe._006_ ;
 wire \AuI.pe._007_ ;
 wire \AuI.pe._008_ ;
 wire \AuI.pe._009_ ;
 wire \AuI.pe._010_ ;
 wire \AuI.pe._011_ ;
 wire \AuI.pe._012_ ;
 wire \AuI.pe._013_ ;
 wire \AuI.pe._014_ ;
 wire \AuI.pe._015_ ;
 wire \AuI.pe._016_ ;
 wire \AuI.pe._017_ ;
 wire \AuI.pe._018_ ;
 wire \AuI.pe._019_ ;
 wire \AuI.pe._020_ ;
 wire \AuI.pe._021_ ;
 wire \AuI.pe._022_ ;
 wire \AuI.pe._023_ ;
 wire \AuI.pe._024_ ;
 wire \AuI.pe._025_ ;
 wire \AuI.pe._026_ ;
 wire \AuI.pe._027_ ;
 wire \AuI.pe._028_ ;
 wire \AuI.pe._029_ ;
 wire \AuI.pe._030_ ;
 wire \AuI.pe._031_ ;
 wire \AuI.pe._032_ ;
 wire \AuI.pe._033_ ;
 wire \AuI.pe._034_ ;
 wire \AuI.pe._035_ ;
 wire \AuI.pe._036_ ;
 wire \AuI.pe._037_ ;
 wire \AuI.pe._038_ ;
 wire \AuI.pe._039_ ;
 wire \AuI.pe._040_ ;
 wire \AuI.pe._041_ ;
 wire \AuI.pe._042_ ;
 wire \AuI.pe._043_ ;
 wire \AuI.pe._044_ ;
 wire \AuI.pe._045_ ;
 wire \AuI.pe._046_ ;
 wire \AuI.pe._047_ ;
 wire \AuI.pe._048_ ;
 wire \AuI.pe._049_ ;
 wire \AuI.pe._050_ ;
 wire \AuI.pe._051_ ;
 wire \AuI.pe._052_ ;
 wire \AuI.pe._053_ ;
 wire \AuI.pe._054_ ;
 wire \AuI.pe._055_ ;
 wire \AuI.pe._056_ ;
 wire \AuI.pe._057_ ;
 wire \AuI.pe._058_ ;
 wire \AuI.pe._059_ ;
 wire \AuI.pe._060_ ;
 wire \AuI.pe._061_ ;
 wire \AuI.pe._062_ ;
 wire \AuI.pe._063_ ;
 wire \AuI.pe._064_ ;
 wire \AuI.pe._065_ ;
 wire \AuI.pe._066_ ;
 wire \AuI.pe._067_ ;
 wire \AuI.pe._068_ ;
 wire \AuI.pe._069_ ;
 wire \AuI.pe._070_ ;
 wire \AuI.pe._071_ ;
 wire \AuI.pe._072_ ;
 wire \AuI.pe._073_ ;
 wire \AuI.pe._074_ ;
 wire \AuI.pe._075_ ;
 wire \AuI.pe._076_ ;
 wire \AuI.pe._077_ ;
 wire \AuI.pe._078_ ;
 wire \AuI.pe._079_ ;
 wire \AuI.pe._080_ ;
 wire \AuI.pe._081_ ;
 wire \AuI.pe._082_ ;
 wire \AuI.pe._083_ ;
 wire \AuI.pe._084_ ;
 wire \AuI.pe._085_ ;
 wire \AuI.pe._086_ ;
 wire \AuI.pe._087_ ;
 wire \AuI.pe._088_ ;
 wire \AuI.pe._089_ ;
 wire \AuI.pe._090_ ;
 wire \AuI.pe._091_ ;
 wire \AuI.pe._092_ ;
 wire \AuI.pe._093_ ;
 wire \AuI.pe._094_ ;
 wire \AuI.pe._095_ ;
 wire \AuI.pe._096_ ;
 wire \AuI.pe._097_ ;
 wire \AuI.pe._098_ ;
 wire \AuI.pe._099_ ;
 wire \AuI.pe._100_ ;
 wire \AuI.pe._101_ ;
 wire \AuI.pe._102_ ;
 wire \AuI.pe._103_ ;
 wire \AuI.pe._104_ ;
 wire \AuI.pe._105_ ;
 wire \AuI.pe._106_ ;
 wire \AuI.pe._107_ ;
 wire \AuI.pe._108_ ;
 wire \AuI.pe._109_ ;
 wire \AuI.pe._110_ ;
 wire \AuI.pe._111_ ;
 wire \AuI.pe._112_ ;
 wire \AuI.pe._113_ ;
 wire \AuI.pe._114_ ;
 wire \AuI.pe._115_ ;
 wire \AuI.pe._116_ ;
 wire \AuI.pe._117_ ;
 wire \AuI.pe._118_ ;
 wire \AuI.pe._119_ ;
 wire \AuI.pe._120_ ;
 wire \AuI.pe._121_ ;
 wire \AuI.pe._122_ ;
 wire \AuI.pe._123_ ;
 wire \AuI.pe._124_ ;
 wire \AuI.pe._125_ ;
 wire \AuI.pe._126_ ;
 wire \AuI.pe._127_ ;
 wire \AuI.pe._128_ ;
 wire \AuI.pe._129_ ;
 wire \AuI.pe._130_ ;
 wire \AuI.pe._131_ ;
 wire \AuI.pe._132_ ;
 wire \AuI.pe._133_ ;
 wire \AuI.pe._134_ ;
 wire \AuI.pe._135_ ;
 wire \AuI.pe._136_ ;
 wire \AuI.pe._137_ ;
 wire \AuI.pe._138_ ;
 wire \AuI.pe._139_ ;
 wire \AuI.pe._140_ ;
 wire \AuI.pe._141_ ;
 wire \AuI.pe._142_ ;
 wire \AuI.pe._143_ ;
 wire \AuI.pe._144_ ;
 wire \AuI.pe._145_ ;
 wire \AuI.pe._146_ ;
 wire \AuI.pe._147_ ;
 wire \AuI.pe._148_ ;
 wire \AuI.pe._149_ ;
 wire \AuI.pe._150_ ;
 wire \AuI.pe._151_ ;
 wire \AuI.pe._152_ ;
 wire \AuI.pe._153_ ;
 wire \AuI.pe._154_ ;
 wire \AuI.pe._155_ ;
 wire \AuI.pe._156_ ;
 wire \AuI.pe._157_ ;
 wire \AuI.pe._158_ ;
 wire \AuI.pe._159_ ;
 wire \AuI.pe._160_ ;
 wire \AuI.pe._161_ ;
 wire \AuI.pe._162_ ;
 wire \AuI.pe._163_ ;
 wire \AuI.pe._164_ ;
 wire \AuI.pe._165_ ;
 wire \AuI.pe._166_ ;
 wire \AuI.pe._167_ ;
 wire \AuI.pe._168_ ;
 wire \AuI.pe._169_ ;
 wire \AuI.pe._170_ ;
 wire \AuI.pe._171_ ;
 wire \AuI.pe._172_ ;
 wire \AuI.pe._173_ ;
 wire \AuI.pe._174_ ;
 wire \AuI.pe._175_ ;
 wire \AuI.pe._176_ ;
 wire \AuI.pe._177_ ;
 wire \AuI.pe._178_ ;
 wire \AuI.pe._179_ ;
 wire \AuI.pe._180_ ;
 wire \AuI.pe._181_ ;
 wire \AuI.pe._182_ ;
 wire \AuI.pe._183_ ;
 wire \AuI.pe._184_ ;
 wire \AuI.pe._185_ ;
 wire \AuI.pe._186_ ;
 wire \AuI.pe._187_ ;
 wire \AuI.pe._188_ ;
 wire \AuI.pe._189_ ;
 wire \AuI.pe._190_ ;
 wire \AuI.pe._191_ ;
 wire \AuI.pe._192_ ;
 wire \AuI.pe._193_ ;
 wire \AuI.pe._194_ ;
 wire \AuI.pe._195_ ;
 wire \AuI.pe._196_ ;
 wire \AuI.pe._197_ ;
 wire \AuI.pe._198_ ;
 wire \AuI.pe._199_ ;
 wire \AuI.pe._200_ ;
 wire \AuI.pe._201_ ;
 wire \AuI.pe._202_ ;
 wire \AuI.pe._203_ ;
 wire \AuI.pe._204_ ;
 wire \AuI.pe._205_ ;
 wire \AuI.pe._206_ ;
 wire \AuI.pe._207_ ;
 wire \AuI.pe._208_ ;
 wire \AuI.pe._209_ ;
 wire \AuI.pe._210_ ;
 wire \AuI.pe._211_ ;
 wire \AuI.pe._212_ ;
 wire \AuI.pe._213_ ;
 wire \AuI.pe._214_ ;
 wire \AuI.pe._215_ ;
 wire \AuI.pe._216_ ;
 wire \AuI.pe._217_ ;
 wire \AuI.pe._218_ ;
 wire \AuI.pe._219_ ;
 wire \AuI.pe._220_ ;
 wire \AuI.pe._221_ ;
 wire \AuI.pe._222_ ;
 wire \AuI.pe._223_ ;
 wire \AuI.pe._224_ ;
 wire \AuI.pe._225_ ;
 wire \AuI.pe._226_ ;
 wire \AuI.pe._227_ ;
 wire \AuI.pe._228_ ;
 wire \AuI.pe._229_ ;
 wire \AuI.pe._230_ ;
 wire \AuI.pe._231_ ;
 wire \AuI.pe._232_ ;
 wire \AuI.pe._233_ ;
 wire \AuI.pe._234_ ;
 wire \AuI.pe._235_ ;
 wire \AuI.pe._236_ ;
 wire \AuI.pe._237_ ;
 wire \AuI.pe._238_ ;
 wire \AuI.pe._239_ ;
 wire \AuI.pe._240_ ;
 wire \AuI.pe._241_ ;
 wire \AuI.pe._242_ ;
 wire \AuI.pe._243_ ;
 wire \AuI.pe._244_ ;
 wire \AuI.pe._245_ ;
 wire \AuI.pe._246_ ;
 wire \AuI.pe._247_ ;
 wire \AuI.pe._248_ ;
 wire \AuI.pe._249_ ;
 wire \AuI.pe._250_ ;
 wire \AuI.pe._251_ ;
 wire \AuI.pe._252_ ;
 wire \AuI.pe._253_ ;
 wire \AuI.pe._254_ ;
 wire \AuI.pe._255_ ;
 wire \AuI.pe._256_ ;
 wire \AuI.pe._257_ ;
 wire \AuI.pe._258_ ;
 wire \AuI.pe._259_ ;
 wire \AuI.pe._260_ ;
 wire \AuI.pe._261_ ;
 wire \AuI.pe._262_ ;
 wire \AuI.pe._263_ ;
 wire \AuI.pe._264_ ;
 wire \AuI.pe._265_ ;
 wire \AuI.pe._266_ ;
 wire \AuI.pe._267_ ;
 wire \AuI.pe._268_ ;
 wire \AuI.pe._269_ ;
 wire \AuI.pe._270_ ;
 wire \AuI.pe._271_ ;
 wire \AuI.pe._272_ ;
 wire \AuI.pe._273_ ;
 wire \AuI.pe._274_ ;
 wire \AuI.pe._275_ ;
 wire \AuI.pe._276_ ;
 wire \AuI.pe._277_ ;
 wire \AuI.pe._278_ ;
 wire \AuI.pe._279_ ;
 wire \AuI.pe._280_ ;
 wire \AuI.pe._281_ ;
 wire \AuI.pe._282_ ;
 wire \AuI.pe._283_ ;
 wire \AuI.pe._284_ ;
 wire \AuI.pe._285_ ;
 wire \AuI.pe._286_ ;
 wire \AuI.pe._287_ ;
 wire \AuI.pe._288_ ;
 wire \AuI.pe._289_ ;
 wire \AuI.pe._290_ ;
 wire \AuI.pe._291_ ;
 wire \AuI.pe._292_ ;
 wire \AuI.pe._293_ ;
 wire \AuI.pe._294_ ;
 wire \AuI.pe._295_ ;
 wire \AuI.pe._296_ ;
 wire \AuI.pe._297_ ;
 wire \AuI.pe._298_ ;
 wire \AuI.pe._299_ ;
 wire \AuI.pe._300_ ;
 wire \AuI.pe._301_ ;
 wire \AuI.pe._302_ ;
 wire \AuI.pe._303_ ;
 wire \AuI.pe._304_ ;
 wire \AuI.pe._305_ ;
 wire \AuI.pe._306_ ;
 wire \AuI.pe._307_ ;
 wire \AuI.pe._308_ ;
 wire \AuI.pe._309_ ;
 wire \AuI.pe._310_ ;
 wire \AuI.pe._311_ ;
 wire \AuI.pe._312_ ;
 wire \AuI.pe._313_ ;
 wire \AuI.pe._314_ ;
 wire \AuI.pe._318_ ;
 wire \AuI.pe._319_ ;
 wire \AuI.pe._320_ ;
 wire \AuI.pe._321_ ;
 wire \AuI.pe._322_ ;
 wire \AuI.pe._323_ ;
 wire \AuI.pe._324_ ;
 wire \AuI.pe._325_ ;
 wire \AuI.pe._326_ ;
 wire \AuI.pe._327_ ;
 wire \AuI.pe._328_ ;
 wire \AuI.pe._329_ ;
 wire \AuI.pe._330_ ;
 wire \AuI.pe._331_ ;
 wire \AuI.pe._332_ ;
 wire \AuI.pe._333_ ;
 wire \AuI.pe._334_ ;
 wire \AuI.pe._335_ ;
 wire \AuI.pe._336_ ;
 wire \AuI.pe._337_ ;
 wire \AuI.pe._338_ ;
 wire \AuI.pe._339_ ;
 wire \AuI.pe._340_ ;
 wire \AuI.pe._341_ ;
 wire \AuI.pe._342_ ;
 wire \AuI.pe._343_ ;
 wire \AuI.pe._344_ ;
 wire \AuI.pe._345_ ;
 wire \AuI.pe._346_ ;
 wire \AuI.pe._347_ ;
 wire \AuI.pe._348_ ;
 wire \AuI.pe._349_ ;
 wire \AuI.pe._350_ ;
 wire \AuI.pe._351_ ;
 wire \AuI.pe._352_ ;
 wire \AuI.pe._353_ ;
 wire \AuI.pe._354_ ;
 wire \AuI.pe._355_ ;
 wire \AuI.pe._356_ ;
 wire \AuI.pe._357_ ;
 wire \AuI.pe._358_ ;
 wire \AuI.pe._359_ ;
 wire \AuI.pe._360_ ;
 wire \AuI.pe._361_ ;
 wire \AuI.pe._362_ ;
 wire \AuI.pe._363_ ;
 wire \AuI.pe._364_ ;
 wire \AuI.pe._365_ ;
 wire \AuI.pe._366_ ;
 wire \AuI.pe._367_ ;
 wire \AuI.pe._368_ ;
 wire \AuI.pe._369_ ;
 wire \AuI.pe._370_ ;
 wire \AuI.pe._371_ ;
 wire \AuI.pe._372_ ;
 wire \AuI.pe._373_ ;
 wire \AuI.pe._374_ ;
 wire \AuI.pe._375_ ;
 wire \AuI.pe._376_ ;
 wire \AuI.pe._377_ ;
 wire \AuI.pe._378_ ;
 wire \AuI.pe._379_ ;
 wire \AuI.pe._380_ ;
 wire \AuI.pe._381_ ;
 wire \AuI.pe._382_ ;
 wire \AuI.pe._383_ ;
 wire \AuI.pe._384_ ;
 wire \AuI.pe._385_ ;
 wire \AuI.pe._386_ ;
 wire \AuI.pe._387_ ;
 wire \AuI.pe._388_ ;
 wire \AuI.pe._389_ ;
 wire \AuI.pe._390_ ;
 wire \AuI.pe._391_ ;
 wire \AuI.pe._392_ ;
 wire \AuI.pe._393_ ;
 wire \AuI.pe._394_ ;
 wire \AuI.pe._395_ ;
 wire \AuI.pe._396_ ;
 wire \AuI.pe._397_ ;
 wire \AuI.pe._398_ ;
 wire \AuI.pe._399_ ;
 wire \AuI.pe.significand[0] ;
 wire \AuI.pe.significand[10] ;
 wire \AuI.pe.significand[11] ;
 wire \AuI.pe.significand[12] ;
 wire \AuI.pe.significand[13] ;
 wire \AuI.pe.significand[14] ;
 wire \AuI.pe.significand[15] ;
 wire \AuI.pe.significand[16] ;
 wire \AuI.pe.significand[17] ;
 wire \AuI.pe.significand[18] ;
 wire \AuI.pe.significand[19] ;
 wire \AuI.pe.significand[1] ;
 wire \AuI.pe.significand[20] ;
 wire \AuI.pe.significand[21] ;
 wire \AuI.pe.significand[22] ;
 wire \AuI.pe.significand[23] ;
 wire \AuI.pe.significand[24] ;
 wire \AuI.pe.significand[2] ;
 wire \AuI.pe.significand[3] ;
 wire \AuI.pe.significand[4] ;
 wire \AuI.pe.significand[5] ;
 wire \AuI.pe.significand[6] ;
 wire \AuI.pe.significand[7] ;
 wire \AuI.pe.significand[8] ;
 wire \AuI.pe.significand[9] ;
 wire \AuI.result[0] ;
 wire \AuI.result[10] ;
 wire \AuI.result[11] ;
 wire \AuI.result[12] ;
 wire \AuI.result[13] ;
 wire \AuI.result[14] ;
 wire \AuI.result[15] ;
 wire \AuI.result[16] ;
 wire \AuI.result[17] ;
 wire \AuI.result[18] ;
 wire \AuI.result[19] ;
 wire \AuI.result[1] ;
 wire \AuI.result[20] ;
 wire \AuI.result[21] ;
 wire \AuI.result[22] ;
 wire \AuI.result[23] ;
 wire \AuI.result[24] ;
 wire \AuI.result[25] ;
 wire \AuI.result[26] ;
 wire \AuI.result[27] ;
 wire \AuI.result[28] ;
 wire \AuI.result[29] ;
 wire \AuI.result[2] ;
 wire \AuI.result[30] ;
 wire \AuI.result[31] ;
 wire \AuI.result[3] ;
 wire \AuI.result[4] ;
 wire \AuI.result[5] ;
 wire \AuI.result[6] ;
 wire \AuI.result[7] ;
 wire \AuI.result[8] ;
 wire \AuI.result[9] ;
 wire \FuI.Integer[0] ;
 wire \FuI.Integer[10] ;
 wire \FuI.Integer[11] ;
 wire \FuI.Integer[12] ;
 wire \FuI.Integer[13] ;
 wire \FuI.Integer[14] ;
 wire \FuI.Integer[15] ;
 wire \FuI.Integer[16] ;
 wire \FuI.Integer[17] ;
 wire \FuI.Integer[18] ;
 wire \FuI.Integer[19] ;
 wire \FuI.Integer[1] ;
 wire \FuI.Integer[20] ;
 wire \FuI.Integer[21] ;
 wire net135;
 wire \FuI.Integer[23] ;
 wire \FuI.Integer[24] ;
 wire \FuI.Integer[25] ;
 wire \FuI.Integer[26] ;
 wire \FuI.Integer[27] ;
 wire \FuI.Integer[28] ;
 wire \FuI.Integer[29] ;
 wire \FuI.Integer[2] ;
 wire \FuI.Integer[30] ;
 wire \FuI.Integer[31] ;
 wire \FuI.Integer[3] ;
 wire \FuI.Integer[4] ;
 wire \FuI.Integer[5] ;
 wire \FuI.Integer[6] ;
 wire \FuI.Integer[7] ;
 wire \FuI.Integer[8] ;
 wire \FuI.Integer[9] ;
 wire \FuI._000_ ;
 wire \FuI._001_ ;
 wire \FuI._002_ ;
 wire \FuI._003_ ;
 wire \FuI._004_ ;
 wire \FuI._005_ ;
 wire \FuI._006_ ;
 wire \FuI._007_ ;
 wire \FuI._008_ ;
 wire \FuI._009_ ;
 wire \FuI._010_ ;
 wire \FuI._011_ ;
 wire \FuI._012_ ;
 wire \FuI._013_ ;
 wire \FuI._014_ ;
 wire \FuI._015_ ;
 wire \FuI._016_ ;
 wire \FuI._017_ ;
 wire \FuI._018_ ;
 wire \FuI._019_ ;
 wire \FuI._020_ ;
 wire \FuI._021_ ;
 wire \FuI._023_ ;
 wire \FuI._024_ ;
 wire \FuI._025_ ;
 wire \FuI._026_ ;
 wire \FuI._027_ ;
 wire \FuI._028_ ;
 wire \FuI._029_ ;
 wire \FuI._030_ ;
 wire \FuI._031_ ;
 wire \FuI._032_ ;
 wire \FuI._033_ ;
 wire \FuI._034_ ;
 wire \FuI._035_ ;
 wire \FuI._036_ ;
 wire \FuI._037_ ;
 wire \FuI._038_ ;
 wire \FuI._039_ ;
 wire \FuI._040_ ;
 wire \FuI._041_ ;
 wire \FuI._042_ ;
 wire \FuI._043_ ;
 wire \FuI._044_ ;
 wire \FuI._045_ ;
 wire \FuI._046_ ;
 wire \FuI._047_ ;
 wire \FuI._048_ ;
 wire \FuI._049_ ;
 wire \FuI._050_ ;
 wire \FuI._051_ ;
 wire \FuI._052_ ;
 wire \FuI._053_ ;
 wire \FuI._054_ ;
 wire \FuI._055_ ;
 wire \FuI._056_ ;
 wire \FuI._057_ ;
 wire \FuI._058_ ;
 wire \FuI._059_ ;
 wire \FuI._060_ ;
 wire \FuI._061_ ;
 wire \FuI._062_ ;
 wire \FuI._063_ ;
 wire \FuI._064_ ;
 wire \FuI.a_operand[10] ;
 wire \FuI.a_operand[11] ;
 wire \FuI.a_operand[12] ;
 wire \FuI.a_operand[13] ;
 wire \FuI.a_operand[14] ;
 wire \FuI.a_operand[15] ;
 wire \FuI.a_operand[16] ;
 wire \FuI.a_operand[17] ;
 wire \FuI.a_operand[18] ;
 wire \FuI.a_operand[19] ;
 wire \FuI.a_operand[1] ;
 wire \FuI.a_operand[20] ;
 wire \FuI.a_operand[21] ;
 wire \FuI.a_operand[22] ;
 wire \FuI.a_operand[23] ;
 wire \FuI.a_operand[24] ;
 wire \FuI.a_operand[25] ;
 wire \FuI.a_operand[26] ;
 wire \FuI.a_operand[27] ;
 wire \FuI.a_operand[28] ;
 wire \FuI.a_operand[29] ;
 wire \FuI.a_operand[2] ;
 wire \FuI.a_operand[30] ;
 wire \FuI.a_operand[31] ;
 wire \FuI.a_operand[3] ;
 wire \FuI.a_operand[4] ;
 wire \FuI.a_operand[5] ;
 wire \FuI.a_operand[6] ;
 wire \FuI.a_operand[7] ;
 wire \FuI.a_operand[8] ;
 wire \FuI.a_operand[9] ;
 wire \MuI.Exception ;
 wire \MuI.Overflow ;
 wire \MuI.Underflow ;
 wire \MuI._0000_ ;
 wire \MuI._0001_ ;
 wire \MuI._0002_ ;
 wire \MuI._0003_ ;
 wire \MuI._0004_ ;
 wire \MuI._0005_ ;
 wire \MuI._0006_ ;
 wire \MuI._0007_ ;
 wire \MuI._0008_ ;
 wire \MuI._0009_ ;
 wire \MuI._0010_ ;
 wire \MuI._0011_ ;
 wire \MuI._0012_ ;
 wire \MuI._0013_ ;
 wire \MuI._0014_ ;
 wire \MuI._0015_ ;
 wire \MuI._0016_ ;
 wire \MuI._0017_ ;
 wire \MuI._0018_ ;
 wire \MuI._0019_ ;
 wire \MuI._0020_ ;
 wire \MuI._0021_ ;
 wire \MuI._0022_ ;
 wire \MuI._0023_ ;
 wire \MuI._0024_ ;
 wire \MuI._0025_ ;
 wire \MuI._0026_ ;
 wire \MuI._0027_ ;
 wire \MuI._0028_ ;
 wire \MuI._0029_ ;
 wire \MuI._0030_ ;
 wire \MuI._0031_ ;
 wire \MuI._0032_ ;
 wire \MuI._0033_ ;
 wire \MuI._0034_ ;
 wire \MuI._0035_ ;
 wire \MuI._0036_ ;
 wire \MuI._0037_ ;
 wire \MuI._0038_ ;
 wire \MuI._0039_ ;
 wire \MuI._0040_ ;
 wire \MuI._0041_ ;
 wire \MuI._0042_ ;
 wire \MuI._0043_ ;
 wire \MuI._0044_ ;
 wire \MuI._0045_ ;
 wire \MuI._0046_ ;
 wire \MuI._0047_ ;
 wire \MuI._0048_ ;
 wire \MuI._0049_ ;
 wire \MuI._0050_ ;
 wire \MuI._0051_ ;
 wire \MuI._0052_ ;
 wire \MuI._0053_ ;
 wire \MuI._0054_ ;
 wire \MuI._0055_ ;
 wire \MuI._0056_ ;
 wire \MuI._0057_ ;
 wire \MuI._0058_ ;
 wire \MuI._0059_ ;
 wire \MuI._0060_ ;
 wire \MuI._0061_ ;
 wire \MuI._0062_ ;
 wire \MuI._0063_ ;
 wire \MuI._0064_ ;
 wire \MuI._0065_ ;
 wire \MuI._0066_ ;
 wire \MuI._0067_ ;
 wire \MuI._0068_ ;
 wire \MuI._0069_ ;
 wire \MuI._0070_ ;
 wire \MuI._0071_ ;
 wire \MuI._0072_ ;
 wire \MuI._0073_ ;
 wire \MuI._0074_ ;
 wire \MuI._0075_ ;
 wire \MuI._0076_ ;
 wire \MuI._0077_ ;
 wire \MuI._0078_ ;
 wire \MuI._0079_ ;
 wire \MuI._0080_ ;
 wire \MuI._0081_ ;
 wire \MuI._0082_ ;
 wire \MuI._0083_ ;
 wire \MuI._0084_ ;
 wire \MuI._0085_ ;
 wire \MuI._0086_ ;
 wire \MuI._0087_ ;
 wire \MuI._0088_ ;
 wire \MuI._0089_ ;
 wire \MuI._0090_ ;
 wire \MuI._0091_ ;
 wire \MuI._0092_ ;
 wire \MuI._0093_ ;
 wire \MuI._0094_ ;
 wire \MuI._0095_ ;
 wire \MuI._0096_ ;
 wire \MuI._0097_ ;
 wire \MuI._0098_ ;
 wire \MuI._0099_ ;
 wire \MuI._0100_ ;
 wire \MuI._0101_ ;
 wire \MuI._0102_ ;
 wire \MuI._0103_ ;
 wire \MuI._0104_ ;
 wire \MuI._0105_ ;
 wire \MuI._0106_ ;
 wire \MuI._0107_ ;
 wire \MuI._0108_ ;
 wire \MuI._0109_ ;
 wire \MuI._0110_ ;
 wire \MuI._0111_ ;
 wire \MuI._0112_ ;
 wire \MuI._0113_ ;
 wire \MuI._0114_ ;
 wire \MuI._0115_ ;
 wire \MuI._0116_ ;
 wire \MuI._0117_ ;
 wire \MuI._0118_ ;
 wire \MuI._0119_ ;
 wire \MuI._0120_ ;
 wire \MuI._0121_ ;
 wire \MuI._0122_ ;
 wire \MuI._0123_ ;
 wire \MuI._0124_ ;
 wire \MuI._0125_ ;
 wire \MuI._0126_ ;
 wire \MuI._0127_ ;
 wire \MuI._0128_ ;
 wire \MuI._0129_ ;
 wire \MuI._0130_ ;
 wire \MuI._0131_ ;
 wire \MuI._0132_ ;
 wire \MuI._0133_ ;
 wire \MuI._0134_ ;
 wire \MuI._0135_ ;
 wire \MuI._0136_ ;
 wire \MuI._0137_ ;
 wire \MuI._0138_ ;
 wire \MuI._0139_ ;
 wire \MuI._0140_ ;
 wire \MuI._0141_ ;
 wire \MuI._0142_ ;
 wire \MuI._0143_ ;
 wire \MuI._0144_ ;
 wire \MuI._0145_ ;
 wire \MuI._0146_ ;
 wire \MuI._0147_ ;
 wire \MuI._0148_ ;
 wire \MuI._0149_ ;
 wire \MuI._0150_ ;
 wire \MuI._0151_ ;
 wire \MuI._0152_ ;
 wire \MuI._0153_ ;
 wire \MuI._0154_ ;
 wire \MuI._0155_ ;
 wire \MuI._0156_ ;
 wire \MuI._0157_ ;
 wire \MuI._0158_ ;
 wire \MuI._0159_ ;
 wire \MuI._0160_ ;
 wire \MuI._0161_ ;
 wire \MuI._0162_ ;
 wire \MuI._0163_ ;
 wire \MuI._0164_ ;
 wire \MuI._0165_ ;
 wire \MuI._0166_ ;
 wire \MuI._0167_ ;
 wire \MuI._0168_ ;
 wire \MuI._0169_ ;
 wire \MuI._0170_ ;
 wire \MuI._0171_ ;
 wire \MuI._0172_ ;
 wire \MuI._0173_ ;
 wire \MuI._0174_ ;
 wire \MuI._0175_ ;
 wire \MuI._0176_ ;
 wire \MuI._0177_ ;
 wire \MuI._0178_ ;
 wire \MuI._0179_ ;
 wire \MuI._0180_ ;
 wire \MuI._0181_ ;
 wire \MuI._0182_ ;
 wire \MuI._0183_ ;
 wire \MuI._0184_ ;
 wire \MuI._0185_ ;
 wire \MuI._0186_ ;
 wire \MuI._0187_ ;
 wire \MuI._0188_ ;
 wire \MuI._0189_ ;
 wire \MuI._0190_ ;
 wire \MuI._0191_ ;
 wire \MuI._0192_ ;
 wire \MuI._0193_ ;
 wire \MuI._0194_ ;
 wire \MuI._0195_ ;
 wire \MuI._0196_ ;
 wire \MuI._0197_ ;
 wire \MuI._0198_ ;
 wire \MuI._0199_ ;
 wire \MuI._0200_ ;
 wire \MuI._0201_ ;
 wire \MuI._0202_ ;
 wire \MuI._0203_ ;
 wire \MuI._0204_ ;
 wire \MuI._0205_ ;
 wire \MuI._0206_ ;
 wire \MuI._0207_ ;
 wire \MuI._0208_ ;
 wire \MuI._0209_ ;
 wire \MuI._0210_ ;
 wire \MuI._0211_ ;
 wire \MuI._0212_ ;
 wire \MuI._0213_ ;
 wire \MuI._0214_ ;
 wire \MuI._0215_ ;
 wire \MuI._0216_ ;
 wire \MuI._0217_ ;
 wire \MuI._0218_ ;
 wire \MuI._0219_ ;
 wire \MuI._0220_ ;
 wire \MuI._0221_ ;
 wire \MuI._0222_ ;
 wire \MuI._0223_ ;
 wire \MuI._0224_ ;
 wire \MuI._0225_ ;
 wire \MuI._0226_ ;
 wire \MuI._0227_ ;
 wire \MuI._0228_ ;
 wire \MuI._0229_ ;
 wire \MuI._0230_ ;
 wire \MuI._0231_ ;
 wire \MuI._0232_ ;
 wire \MuI._0233_ ;
 wire \MuI._0234_ ;
 wire \MuI._0235_ ;
 wire \MuI._0236_ ;
 wire \MuI._0237_ ;
 wire \MuI._0238_ ;
 wire \MuI._0239_ ;
 wire \MuI._0240_ ;
 wire \MuI._0241_ ;
 wire \MuI._0242_ ;
 wire \MuI._0243_ ;
 wire \MuI._0244_ ;
 wire \MuI._0245_ ;
 wire \MuI._0246_ ;
 wire \MuI._0247_ ;
 wire \MuI._0248_ ;
 wire \MuI._0249_ ;
 wire \MuI._0250_ ;
 wire \MuI._0251_ ;
 wire \MuI._0252_ ;
 wire \MuI._0253_ ;
 wire \MuI._0254_ ;
 wire \MuI._0255_ ;
 wire \MuI._0256_ ;
 wire \MuI._0257_ ;
 wire \MuI._0258_ ;
 wire \MuI._0259_ ;
 wire \MuI._0260_ ;
 wire \MuI._0261_ ;
 wire \MuI._0262_ ;
 wire \MuI._0263_ ;
 wire \MuI._0264_ ;
 wire \MuI._0265_ ;
 wire \MuI._0266_ ;
 wire \MuI._0267_ ;
 wire \MuI._0268_ ;
 wire \MuI._0269_ ;
 wire \MuI._0270_ ;
 wire \MuI._0271_ ;
 wire \MuI._0272_ ;
 wire \MuI._0273_ ;
 wire \MuI._0274_ ;
 wire \MuI._0275_ ;
 wire \MuI._0276_ ;
 wire \MuI._0277_ ;
 wire \MuI._0278_ ;
 wire \MuI._0279_ ;
 wire \MuI._0280_ ;
 wire \MuI._0281_ ;
 wire \MuI._0282_ ;
 wire \MuI._0283_ ;
 wire \MuI._0284_ ;
 wire \MuI._0285_ ;
 wire \MuI._0286_ ;
 wire \MuI._0287_ ;
 wire \MuI._0288_ ;
 wire \MuI._0289_ ;
 wire \MuI._0290_ ;
 wire \MuI._0291_ ;
 wire \MuI._0292_ ;
 wire \MuI._0293_ ;
 wire \MuI._0294_ ;
 wire \MuI._0295_ ;
 wire \MuI._0296_ ;
 wire \MuI._0297_ ;
 wire \MuI._0298_ ;
 wire \MuI._0299_ ;
 wire \MuI._0300_ ;
 wire \MuI._0301_ ;
 wire \MuI._0302_ ;
 wire \MuI._0303_ ;
 wire \MuI._0304_ ;
 wire \MuI._0305_ ;
 wire \MuI._0306_ ;
 wire \MuI._0307_ ;
 wire \MuI._0308_ ;
 wire \MuI._0309_ ;
 wire \MuI._0310_ ;
 wire \MuI._0311_ ;
 wire \MuI._0312_ ;
 wire \MuI._0313_ ;
 wire \MuI._0314_ ;
 wire \MuI._0315_ ;
 wire \MuI._0316_ ;
 wire \MuI._0317_ ;
 wire \MuI._0318_ ;
 wire \MuI._0319_ ;
 wire \MuI._0320_ ;
 wire \MuI._0321_ ;
 wire \MuI._0322_ ;
 wire \MuI._0323_ ;
 wire \MuI._0324_ ;
 wire \MuI._0325_ ;
 wire \MuI._0326_ ;
 wire \MuI._0327_ ;
 wire \MuI._0328_ ;
 wire \MuI._0329_ ;
 wire \MuI._0330_ ;
 wire \MuI._0331_ ;
 wire \MuI._0332_ ;
 wire \MuI._0333_ ;
 wire \MuI._0334_ ;
 wire \MuI._0335_ ;
 wire \MuI._0336_ ;
 wire \MuI._0337_ ;
 wire \MuI._0338_ ;
 wire \MuI._0339_ ;
 wire \MuI._0340_ ;
 wire \MuI._0341_ ;
 wire \MuI._0342_ ;
 wire \MuI._0343_ ;
 wire \MuI._0344_ ;
 wire \MuI._0345_ ;
 wire \MuI._0346_ ;
 wire \MuI._0347_ ;
 wire \MuI._0348_ ;
 wire \MuI._0349_ ;
 wire \MuI._0350_ ;
 wire \MuI._0351_ ;
 wire \MuI._0352_ ;
 wire \MuI._0353_ ;
 wire \MuI._0354_ ;
 wire \MuI._0355_ ;
 wire \MuI._0356_ ;
 wire \MuI._0357_ ;
 wire \MuI._0358_ ;
 wire \MuI._0359_ ;
 wire \MuI._0360_ ;
 wire \MuI._0361_ ;
 wire \MuI._0362_ ;
 wire \MuI._0363_ ;
 wire \MuI._0364_ ;
 wire \MuI._0365_ ;
 wire \MuI._0366_ ;
 wire \MuI._0367_ ;
 wire \MuI._0368_ ;
 wire \MuI._0369_ ;
 wire \MuI._0370_ ;
 wire \MuI._0371_ ;
 wire \MuI._0372_ ;
 wire \MuI._0373_ ;
 wire \MuI._0374_ ;
 wire \MuI._0375_ ;
 wire \MuI._0376_ ;
 wire \MuI._0377_ ;
 wire \MuI._0378_ ;
 wire \MuI._0379_ ;
 wire \MuI._0380_ ;
 wire \MuI._0381_ ;
 wire \MuI._0382_ ;
 wire \MuI._0383_ ;
 wire \MuI._0384_ ;
 wire \MuI._0385_ ;
 wire \MuI._0386_ ;
 wire \MuI._0387_ ;
 wire \MuI._0388_ ;
 wire \MuI._0389_ ;
 wire \MuI._0390_ ;
 wire \MuI._0391_ ;
 wire \MuI._0392_ ;
 wire \MuI._0393_ ;
 wire \MuI._0394_ ;
 wire \MuI._0395_ ;
 wire \MuI._0396_ ;
 wire \MuI._0397_ ;
 wire \MuI._0398_ ;
 wire \MuI._0399_ ;
 wire \MuI._0400_ ;
 wire \MuI._0401_ ;
 wire \MuI._0402_ ;
 wire \MuI._0403_ ;
 wire \MuI._0404_ ;
 wire \MuI._0405_ ;
 wire \MuI._0406_ ;
 wire \MuI._0407_ ;
 wire \MuI._0408_ ;
 wire \MuI._0409_ ;
 wire \MuI._0410_ ;
 wire \MuI._0411_ ;
 wire \MuI._0412_ ;
 wire \MuI._0413_ ;
 wire \MuI._0414_ ;
 wire \MuI._0415_ ;
 wire \MuI._0416_ ;
 wire \MuI._0417_ ;
 wire \MuI._0418_ ;
 wire \MuI._0419_ ;
 wire \MuI._0420_ ;
 wire \MuI._0421_ ;
 wire \MuI._0422_ ;
 wire \MuI._0423_ ;
 wire \MuI._0424_ ;
 wire \MuI._0425_ ;
 wire \MuI._0426_ ;
 wire \MuI._0427_ ;
 wire \MuI._0428_ ;
 wire \MuI._0429_ ;
 wire \MuI._0430_ ;
 wire \MuI._0431_ ;
 wire \MuI._0432_ ;
 wire \MuI._0433_ ;
 wire \MuI._0434_ ;
 wire \MuI._0435_ ;
 wire \MuI._0436_ ;
 wire \MuI._0437_ ;
 wire \MuI._0438_ ;
 wire \MuI._0439_ ;
 wire \MuI._0440_ ;
 wire \MuI._0441_ ;
 wire \MuI._0442_ ;
 wire \MuI._0443_ ;
 wire \MuI._0444_ ;
 wire \MuI._0445_ ;
 wire \MuI._0446_ ;
 wire \MuI._0447_ ;
 wire \MuI._0448_ ;
 wire \MuI._0449_ ;
 wire \MuI._0450_ ;
 wire \MuI._0451_ ;
 wire \MuI._0452_ ;
 wire \MuI._0453_ ;
 wire \MuI._0454_ ;
 wire \MuI._0455_ ;
 wire \MuI._0456_ ;
 wire \MuI._0457_ ;
 wire \MuI._0458_ ;
 wire \MuI._0459_ ;
 wire \MuI._0460_ ;
 wire \MuI._0461_ ;
 wire \MuI._0462_ ;
 wire \MuI._0463_ ;
 wire \MuI._0464_ ;
 wire \MuI._0465_ ;
 wire \MuI._0466_ ;
 wire \MuI._0467_ ;
 wire \MuI._0468_ ;
 wire \MuI._0469_ ;
 wire \MuI._0470_ ;
 wire \MuI._0471_ ;
 wire \MuI._0472_ ;
 wire \MuI._0473_ ;
 wire \MuI._0474_ ;
 wire \MuI._0475_ ;
 wire \MuI._0476_ ;
 wire \MuI._0477_ ;
 wire \MuI._0478_ ;
 wire \MuI._0479_ ;
 wire \MuI._0480_ ;
 wire \MuI._0481_ ;
 wire \MuI._0482_ ;
 wire \MuI._0483_ ;
 wire \MuI._0484_ ;
 wire \MuI._0485_ ;
 wire \MuI._0486_ ;
 wire \MuI._0487_ ;
 wire \MuI._0488_ ;
 wire \MuI._0489_ ;
 wire \MuI._0490_ ;
 wire \MuI._0491_ ;
 wire \MuI._0492_ ;
 wire \MuI._0493_ ;
 wire \MuI._0494_ ;
 wire \MuI._0495_ ;
 wire \MuI._0496_ ;
 wire \MuI._0497_ ;
 wire \MuI._0498_ ;
 wire \MuI._0499_ ;
 wire \MuI._0500_ ;
 wire \MuI._0501_ ;
 wire \MuI._0502_ ;
 wire \MuI._0503_ ;
 wire \MuI._0504_ ;
 wire \MuI._0505_ ;
 wire \MuI._0506_ ;
 wire \MuI._0507_ ;
 wire \MuI._0508_ ;
 wire \MuI._0509_ ;
 wire \MuI._0510_ ;
 wire \MuI._0511_ ;
 wire \MuI._0512_ ;
 wire \MuI._0513_ ;
 wire \MuI._0514_ ;
 wire \MuI._0515_ ;
 wire \MuI._0516_ ;
 wire \MuI._0517_ ;
 wire \MuI._0518_ ;
 wire \MuI._0519_ ;
 wire \MuI._0520_ ;
 wire \MuI._0521_ ;
 wire \MuI._0522_ ;
 wire \MuI._0523_ ;
 wire \MuI._0524_ ;
 wire \MuI._0525_ ;
 wire \MuI._0526_ ;
 wire \MuI._0527_ ;
 wire \MuI._0528_ ;
 wire \MuI._0529_ ;
 wire \MuI._0530_ ;
 wire \MuI._0531_ ;
 wire \MuI._0532_ ;
 wire \MuI._0533_ ;
 wire \MuI._0534_ ;
 wire \MuI._0535_ ;
 wire \MuI._0536_ ;
 wire \MuI._0537_ ;
 wire \MuI._0538_ ;
 wire \MuI._0539_ ;
 wire \MuI._0540_ ;
 wire \MuI._0541_ ;
 wire \MuI._0542_ ;
 wire \MuI._0543_ ;
 wire \MuI._0544_ ;
 wire \MuI._0545_ ;
 wire \MuI._0546_ ;
 wire \MuI._0547_ ;
 wire \MuI._0548_ ;
 wire \MuI._0549_ ;
 wire \MuI._0550_ ;
 wire \MuI._0551_ ;
 wire \MuI._0552_ ;
 wire \MuI._0553_ ;
 wire \MuI._0554_ ;
 wire \MuI._0555_ ;
 wire \MuI._0556_ ;
 wire \MuI._0557_ ;
 wire \MuI._0558_ ;
 wire \MuI._0559_ ;
 wire \MuI._0560_ ;
 wire \MuI._0561_ ;
 wire \MuI._0562_ ;
 wire \MuI._0563_ ;
 wire \MuI._0564_ ;
 wire \MuI._0565_ ;
 wire \MuI._0566_ ;
 wire \MuI._0567_ ;
 wire \MuI._0568_ ;
 wire \MuI._0569_ ;
 wire \MuI._0570_ ;
 wire \MuI._0571_ ;
 wire \MuI._0572_ ;
 wire \MuI._0573_ ;
 wire \MuI._0574_ ;
 wire \MuI._0575_ ;
 wire \MuI._0576_ ;
 wire \MuI._0577_ ;
 wire \MuI._0578_ ;
 wire \MuI._0579_ ;
 wire \MuI._0580_ ;
 wire \MuI._0581_ ;
 wire \MuI._0582_ ;
 wire \MuI._0583_ ;
 wire \MuI._0584_ ;
 wire \MuI._0585_ ;
 wire \MuI._0586_ ;
 wire \MuI._0587_ ;
 wire \MuI._0588_ ;
 wire \MuI._0589_ ;
 wire \MuI._0590_ ;
 wire \MuI._0591_ ;
 wire \MuI._0592_ ;
 wire \MuI._0593_ ;
 wire \MuI._0594_ ;
 wire \MuI._0595_ ;
 wire \MuI._0596_ ;
 wire \MuI._0597_ ;
 wire \MuI._0598_ ;
 wire \MuI._0599_ ;
 wire \MuI._0600_ ;
 wire \MuI._0601_ ;
 wire \MuI._0602_ ;
 wire \MuI._0603_ ;
 wire \MuI._0604_ ;
 wire \MuI._0605_ ;
 wire \MuI._0606_ ;
 wire \MuI._0607_ ;
 wire \MuI._0608_ ;
 wire \MuI._0609_ ;
 wire \MuI._0610_ ;
 wire \MuI._0611_ ;
 wire \MuI._0612_ ;
 wire \MuI._0613_ ;
 wire \MuI._0614_ ;
 wire \MuI._0615_ ;
 wire \MuI._0616_ ;
 wire \MuI._0617_ ;
 wire \MuI._0618_ ;
 wire \MuI._0619_ ;
 wire \MuI._0620_ ;
 wire \MuI._0621_ ;
 wire \MuI._0622_ ;
 wire \MuI._0623_ ;
 wire \MuI._0624_ ;
 wire \MuI._0625_ ;
 wire \MuI._0626_ ;
 wire \MuI._0627_ ;
 wire \MuI._0628_ ;
 wire \MuI._0629_ ;
 wire \MuI._0630_ ;
 wire \MuI._0631_ ;
 wire \MuI._0632_ ;
 wire \MuI._0633_ ;
 wire \MuI._0634_ ;
 wire \MuI._0635_ ;
 wire \MuI._0636_ ;
 wire \MuI._0637_ ;
 wire \MuI._0638_ ;
 wire \MuI._0639_ ;
 wire \MuI._0640_ ;
 wire \MuI._0641_ ;
 wire \MuI._0642_ ;
 wire \MuI._0643_ ;
 wire \MuI._0644_ ;
 wire \MuI._0645_ ;
 wire \MuI._0646_ ;
 wire \MuI._0647_ ;
 wire \MuI._0648_ ;
 wire \MuI._0649_ ;
 wire \MuI._0650_ ;
 wire \MuI._0651_ ;
 wire \MuI._0652_ ;
 wire \MuI._0653_ ;
 wire \MuI._0654_ ;
 wire \MuI._0655_ ;
 wire \MuI._0656_ ;
 wire \MuI._0657_ ;
 wire \MuI._0658_ ;
 wire \MuI._0659_ ;
 wire \MuI._0660_ ;
 wire \MuI._0661_ ;
 wire \MuI._0662_ ;
 wire \MuI._0663_ ;
 wire \MuI._0664_ ;
 wire \MuI._0665_ ;
 wire \MuI._0666_ ;
 wire \MuI._0667_ ;
 wire \MuI._0668_ ;
 wire \MuI._0669_ ;
 wire \MuI._0670_ ;
 wire \MuI._0671_ ;
 wire \MuI._0672_ ;
 wire \MuI._0673_ ;
 wire \MuI._0674_ ;
 wire \MuI._0675_ ;
 wire \MuI._0676_ ;
 wire \MuI._0677_ ;
 wire \MuI._0678_ ;
 wire \MuI._0679_ ;
 wire \MuI._0680_ ;
 wire \MuI._0681_ ;
 wire \MuI._0682_ ;
 wire \MuI._0683_ ;
 wire \MuI._0684_ ;
 wire \MuI._0685_ ;
 wire \MuI._0686_ ;
 wire \MuI._0687_ ;
 wire \MuI._0688_ ;
 wire \MuI._0689_ ;
 wire \MuI._0690_ ;
 wire \MuI._0691_ ;
 wire \MuI._0692_ ;
 wire \MuI._0693_ ;
 wire \MuI._0694_ ;
 wire \MuI._0695_ ;
 wire \MuI._0696_ ;
 wire \MuI._0697_ ;
 wire \MuI._0698_ ;
 wire \MuI._0699_ ;
 wire \MuI._0700_ ;
 wire \MuI._0701_ ;
 wire \MuI._0702_ ;
 wire \MuI._0703_ ;
 wire \MuI._0704_ ;
 wire \MuI._0705_ ;
 wire \MuI._0706_ ;
 wire \MuI._0707_ ;
 wire \MuI._0708_ ;
 wire \MuI._0709_ ;
 wire \MuI._0710_ ;
 wire \MuI._0711_ ;
 wire \MuI._0712_ ;
 wire \MuI._0713_ ;
 wire \MuI._0714_ ;
 wire \MuI._0715_ ;
 wire \MuI._0716_ ;
 wire \MuI._0717_ ;
 wire \MuI._0718_ ;
 wire \MuI._0719_ ;
 wire \MuI._0720_ ;
 wire \MuI._0721_ ;
 wire \MuI._0722_ ;
 wire \MuI._0723_ ;
 wire \MuI._0724_ ;
 wire \MuI._0725_ ;
 wire \MuI._0726_ ;
 wire \MuI._0727_ ;
 wire \MuI._0728_ ;
 wire \MuI._0729_ ;
 wire \MuI._0730_ ;
 wire \MuI._0731_ ;
 wire \MuI._0732_ ;
 wire \MuI._0733_ ;
 wire \MuI._0734_ ;
 wire \MuI._0735_ ;
 wire \MuI._0736_ ;
 wire \MuI._0737_ ;
 wire \MuI._0738_ ;
 wire \MuI._0739_ ;
 wire \MuI._0740_ ;
 wire \MuI._0741_ ;
 wire \MuI._0742_ ;
 wire \MuI._0743_ ;
 wire \MuI._0744_ ;
 wire \MuI._0745_ ;
 wire \MuI._0746_ ;
 wire \MuI._0747_ ;
 wire \MuI._0748_ ;
 wire \MuI._0749_ ;
 wire \MuI._0750_ ;
 wire \MuI._0751_ ;
 wire \MuI._0752_ ;
 wire \MuI._0753_ ;
 wire \MuI._0754_ ;
 wire \MuI._0755_ ;
 wire \MuI._0756_ ;
 wire \MuI._0757_ ;
 wire \MuI._0758_ ;
 wire \MuI._0759_ ;
 wire \MuI._0760_ ;
 wire \MuI._0761_ ;
 wire \MuI._0762_ ;
 wire \MuI._0763_ ;
 wire \MuI._0764_ ;
 wire \MuI._0765_ ;
 wire \MuI._0766_ ;
 wire \MuI._0767_ ;
 wire \MuI._0768_ ;
 wire \MuI._0769_ ;
 wire \MuI._0770_ ;
 wire \MuI._0771_ ;
 wire \MuI._0772_ ;
 wire \MuI._0773_ ;
 wire \MuI._0774_ ;
 wire \MuI._0775_ ;
 wire \MuI._0776_ ;
 wire \MuI._0777_ ;
 wire \MuI._0778_ ;
 wire \MuI._0779_ ;
 wire \MuI._0780_ ;
 wire \MuI._0781_ ;
 wire \MuI._0782_ ;
 wire \MuI._0783_ ;
 wire \MuI._0784_ ;
 wire \MuI._0785_ ;
 wire \MuI._0786_ ;
 wire \MuI._0787_ ;
 wire \MuI._0788_ ;
 wire \MuI._0789_ ;
 wire \MuI._0790_ ;
 wire \MuI._0791_ ;
 wire \MuI._0792_ ;
 wire \MuI._0793_ ;
 wire \MuI._0794_ ;
 wire \MuI._0795_ ;
 wire \MuI._0796_ ;
 wire \MuI._0797_ ;
 wire \MuI._0798_ ;
 wire \MuI._0799_ ;
 wire \MuI._0800_ ;
 wire \MuI._0801_ ;
 wire \MuI._0802_ ;
 wire \MuI._0803_ ;
 wire \MuI._0804_ ;
 wire \MuI._0805_ ;
 wire \MuI._0806_ ;
 wire \MuI._0807_ ;
 wire \MuI._0808_ ;
 wire \MuI._0809_ ;
 wire \MuI._0810_ ;
 wire \MuI._0811_ ;
 wire \MuI._0812_ ;
 wire \MuI._0813_ ;
 wire \MuI._0814_ ;
 wire \MuI._0815_ ;
 wire \MuI._0816_ ;
 wire \MuI._0817_ ;
 wire \MuI._0818_ ;
 wire \MuI._0819_ ;
 wire \MuI._0820_ ;
 wire \MuI._0821_ ;
 wire \MuI._0822_ ;
 wire \MuI._0823_ ;
 wire \MuI._0824_ ;
 wire \MuI._0825_ ;
 wire \MuI._0826_ ;
 wire \MuI._0827_ ;
 wire \MuI._0828_ ;
 wire \MuI._0829_ ;
 wire \MuI._0830_ ;
 wire \MuI._0831_ ;
 wire \MuI._0832_ ;
 wire \MuI._0833_ ;
 wire \MuI._0834_ ;
 wire \MuI._0835_ ;
 wire \MuI._0836_ ;
 wire \MuI._0837_ ;
 wire \MuI._0838_ ;
 wire \MuI._0839_ ;
 wire \MuI._0840_ ;
 wire \MuI._0841_ ;
 wire \MuI._0842_ ;
 wire \MuI._0843_ ;
 wire \MuI._0844_ ;
 wire \MuI._0845_ ;
 wire \MuI._0846_ ;
 wire \MuI._0847_ ;
 wire \MuI._0848_ ;
 wire \MuI._0849_ ;
 wire \MuI._0850_ ;
 wire \MuI._0851_ ;
 wire \MuI._0852_ ;
 wire \MuI._0853_ ;
 wire \MuI._0854_ ;
 wire \MuI._0855_ ;
 wire \MuI._0856_ ;
 wire \MuI._0857_ ;
 wire \MuI._0858_ ;
 wire \MuI._0859_ ;
 wire \MuI._0860_ ;
 wire \MuI._0861_ ;
 wire \MuI._0862_ ;
 wire \MuI._0863_ ;
 wire \MuI._0864_ ;
 wire \MuI._0865_ ;
 wire \MuI._0866_ ;
 wire \MuI._0867_ ;
 wire \MuI._0868_ ;
 wire \MuI._0869_ ;
 wire \MuI._0870_ ;
 wire \MuI._0871_ ;
 wire \MuI._0872_ ;
 wire \MuI._0873_ ;
 wire \MuI._0874_ ;
 wire \MuI._0875_ ;
 wire \MuI._0876_ ;
 wire \MuI._0877_ ;
 wire \MuI._0878_ ;
 wire \MuI._0879_ ;
 wire \MuI._0880_ ;
 wire \MuI._0881_ ;
 wire \MuI._0882_ ;
 wire \MuI._0883_ ;
 wire \MuI._0884_ ;
 wire \MuI._0885_ ;
 wire \MuI._0886_ ;
 wire \MuI._0887_ ;
 wire \MuI._0888_ ;
 wire \MuI._0889_ ;
 wire \MuI._0890_ ;
 wire \MuI._0891_ ;
 wire \MuI._0892_ ;
 wire \MuI._0893_ ;
 wire \MuI._0894_ ;
 wire \MuI._0895_ ;
 wire \MuI._0896_ ;
 wire \MuI._0897_ ;
 wire \MuI._0898_ ;
 wire \MuI._0899_ ;
 wire \MuI._0900_ ;
 wire \MuI._0901_ ;
 wire \MuI._0902_ ;
 wire \MuI._0903_ ;
 wire \MuI._0904_ ;
 wire \MuI._0905_ ;
 wire \MuI._0906_ ;
 wire \MuI._0907_ ;
 wire \MuI._0908_ ;
 wire \MuI._0909_ ;
 wire \MuI._0910_ ;
 wire \MuI._0911_ ;
 wire \MuI._0912_ ;
 wire \MuI._0913_ ;
 wire \MuI._0914_ ;
 wire \MuI._0915_ ;
 wire \MuI._0916_ ;
 wire \MuI._0917_ ;
 wire \MuI._0918_ ;
 wire \MuI._0919_ ;
 wire \MuI._0920_ ;
 wire \MuI._0921_ ;
 wire \MuI._0922_ ;
 wire \MuI._0923_ ;
 wire \MuI._0924_ ;
 wire \MuI._0925_ ;
 wire \MuI._0926_ ;
 wire \MuI._0927_ ;
 wire \MuI._0928_ ;
 wire \MuI._0929_ ;
 wire \MuI._0930_ ;
 wire \MuI._0931_ ;
 wire \MuI._0932_ ;
 wire \MuI._0933_ ;
 wire \MuI._0934_ ;
 wire \MuI._0935_ ;
 wire \MuI._0936_ ;
 wire \MuI._0937_ ;
 wire \MuI._0938_ ;
 wire \MuI._0939_ ;
 wire \MuI._0940_ ;
 wire \MuI._0941_ ;
 wire \MuI._0942_ ;
 wire \MuI._0943_ ;
 wire \MuI._0944_ ;
 wire \MuI._0945_ ;
 wire \MuI._0946_ ;
 wire \MuI._0947_ ;
 wire \MuI._0948_ ;
 wire \MuI._0949_ ;
 wire \MuI._0950_ ;
 wire \MuI._0951_ ;
 wire \MuI._0952_ ;
 wire \MuI._0953_ ;
 wire \MuI._0954_ ;
 wire \MuI._0955_ ;
 wire \MuI._0956_ ;
 wire \MuI._0957_ ;
 wire \MuI._0958_ ;
 wire \MuI._0959_ ;
 wire \MuI._0960_ ;
 wire \MuI._0961_ ;
 wire \MuI._0962_ ;
 wire \MuI._0963_ ;
 wire \MuI._0964_ ;
 wire \MuI._0965_ ;
 wire \MuI._0966_ ;
 wire \MuI._0967_ ;
 wire \MuI._0968_ ;
 wire \MuI._0969_ ;
 wire \MuI._0970_ ;
 wire \MuI._0971_ ;
 wire \MuI._0972_ ;
 wire \MuI._0973_ ;
 wire \MuI._0974_ ;
 wire \MuI._0975_ ;
 wire \MuI._0976_ ;
 wire \MuI._0977_ ;
 wire \MuI._0978_ ;
 wire \MuI._0979_ ;
 wire \MuI._0980_ ;
 wire \MuI._0981_ ;
 wire \MuI._0982_ ;
 wire \MuI._0983_ ;
 wire \MuI._0984_ ;
 wire \MuI._0985_ ;
 wire \MuI._0986_ ;
 wire \MuI._0987_ ;
 wire \MuI._0988_ ;
 wire \MuI._0989_ ;
 wire \MuI._0990_ ;
 wire \MuI._0991_ ;
 wire \MuI._0992_ ;
 wire \MuI._0993_ ;
 wire \MuI._0994_ ;
 wire \MuI._0995_ ;
 wire \MuI._0996_ ;
 wire \MuI._0997_ ;
 wire \MuI._0998_ ;
 wire \MuI._0999_ ;
 wire \MuI._1000_ ;
 wire \MuI._1001_ ;
 wire \MuI._1002_ ;
 wire \MuI._1003_ ;
 wire \MuI._1004_ ;
 wire \MuI._1005_ ;
 wire \MuI._1006_ ;
 wire \MuI._1007_ ;
 wire \MuI._1008_ ;
 wire \MuI._1009_ ;
 wire \MuI._1010_ ;
 wire \MuI._1011_ ;
 wire \MuI._1012_ ;
 wire \MuI._1013_ ;
 wire \MuI._1014_ ;
 wire \MuI._1015_ ;
 wire \MuI._1016_ ;
 wire \MuI._1017_ ;
 wire \MuI._1018_ ;
 wire \MuI._1019_ ;
 wire \MuI._1020_ ;
 wire \MuI._1021_ ;
 wire \MuI._1022_ ;
 wire \MuI._1023_ ;
 wire \MuI._1024_ ;
 wire \MuI._1025_ ;
 wire \MuI._1026_ ;
 wire \MuI._1027_ ;
 wire \MuI._1028_ ;
 wire \MuI._1029_ ;
 wire \MuI._1030_ ;
 wire \MuI._1031_ ;
 wire \MuI._1032_ ;
 wire \MuI._1033_ ;
 wire \MuI._1034_ ;
 wire \MuI._1035_ ;
 wire \MuI._1036_ ;
 wire \MuI._1037_ ;
 wire \MuI._1038_ ;
 wire \MuI._1039_ ;
 wire \MuI._1040_ ;
 wire \MuI._1041_ ;
 wire \MuI._1042_ ;
 wire \MuI._1043_ ;
 wire \MuI._1044_ ;
 wire \MuI._1045_ ;
 wire \MuI._1046_ ;
 wire \MuI._1047_ ;
 wire \MuI._1048_ ;
 wire \MuI._1049_ ;
 wire \MuI._1050_ ;
 wire \MuI._1051_ ;
 wire \MuI._1052_ ;
 wire \MuI._1053_ ;
 wire \MuI._1054_ ;
 wire \MuI._1055_ ;
 wire \MuI._1056_ ;
 wire \MuI._1057_ ;
 wire \MuI._1058_ ;
 wire \MuI._1059_ ;
 wire \MuI._1060_ ;
 wire \MuI._1061_ ;
 wire \MuI._1062_ ;
 wire \MuI._1063_ ;
 wire \MuI._1064_ ;
 wire \MuI._1065_ ;
 wire \MuI._1066_ ;
 wire \MuI._1067_ ;
 wire \MuI._1068_ ;
 wire \MuI._1069_ ;
 wire \MuI._1070_ ;
 wire \MuI._1071_ ;
 wire \MuI._1072_ ;
 wire \MuI._1073_ ;
 wire \MuI._1074_ ;
 wire \MuI._1075_ ;
 wire \MuI._1076_ ;
 wire \MuI._1077_ ;
 wire \MuI._1078_ ;
 wire \MuI._1079_ ;
 wire \MuI._1080_ ;
 wire \MuI._1081_ ;
 wire \MuI._1082_ ;
 wire \MuI._1083_ ;
 wire \MuI._1084_ ;
 wire \MuI._1085_ ;
 wire \MuI._1086_ ;
 wire \MuI._1087_ ;
 wire \MuI._1088_ ;
 wire \MuI._1089_ ;
 wire \MuI._1090_ ;
 wire \MuI._1091_ ;
 wire \MuI._1092_ ;
 wire \MuI._1093_ ;
 wire \MuI._1094_ ;
 wire \MuI._1095_ ;
 wire \MuI._1096_ ;
 wire \MuI._1097_ ;
 wire \MuI._1098_ ;
 wire \MuI._1099_ ;
 wire \MuI._1100_ ;
 wire \MuI._1101_ ;
 wire \MuI._1102_ ;
 wire \MuI._1103_ ;
 wire \MuI._1104_ ;
 wire \MuI._1105_ ;
 wire \MuI._1106_ ;
 wire \MuI._1107_ ;
 wire \MuI._1108_ ;
 wire \MuI._1109_ ;
 wire \MuI._1110_ ;
 wire \MuI._1111_ ;
 wire \MuI._1112_ ;
 wire \MuI._1113_ ;
 wire \MuI._1114_ ;
 wire \MuI._1115_ ;
 wire \MuI._1116_ ;
 wire \MuI._1117_ ;
 wire \MuI._1118_ ;
 wire \MuI._1119_ ;
 wire \MuI._1120_ ;
 wire \MuI._1121_ ;
 wire \MuI._1122_ ;
 wire \MuI._1123_ ;
 wire \MuI._1124_ ;
 wire \MuI._1125_ ;
 wire \MuI._1126_ ;
 wire \MuI._1127_ ;
 wire \MuI._1128_ ;
 wire \MuI._1129_ ;
 wire \MuI._1130_ ;
 wire \MuI._1131_ ;
 wire \MuI._1132_ ;
 wire \MuI._1133_ ;
 wire \MuI._1134_ ;
 wire \MuI._1135_ ;
 wire \MuI._1136_ ;
 wire \MuI._1137_ ;
 wire \MuI._1138_ ;
 wire \MuI._1139_ ;
 wire \MuI._1140_ ;
 wire \MuI._1141_ ;
 wire \MuI._1142_ ;
 wire \MuI._1143_ ;
 wire \MuI._1144_ ;
 wire \MuI._1145_ ;
 wire \MuI._1146_ ;
 wire \MuI._1147_ ;
 wire \MuI._1148_ ;
 wire \MuI._1149_ ;
 wire \MuI._1150_ ;
 wire \MuI._1151_ ;
 wire \MuI._1152_ ;
 wire \MuI._1153_ ;
 wire \MuI._1154_ ;
 wire \MuI._1155_ ;
 wire \MuI._1156_ ;
 wire \MuI._1157_ ;
 wire \MuI._1158_ ;
 wire \MuI._1159_ ;
 wire \MuI._1160_ ;
 wire \MuI._1161_ ;
 wire \MuI._1162_ ;
 wire \MuI._1163_ ;
 wire \MuI._1164_ ;
 wire \MuI._1165_ ;
 wire \MuI._1166_ ;
 wire \MuI._1167_ ;
 wire \MuI._1168_ ;
 wire \MuI._1169_ ;
 wire \MuI._1170_ ;
 wire \MuI._1171_ ;
 wire \MuI._1172_ ;
 wire \MuI._1173_ ;
 wire \MuI._1174_ ;
 wire \MuI._1175_ ;
 wire \MuI._1176_ ;
 wire \MuI._1177_ ;
 wire \MuI._1178_ ;
 wire \MuI._1179_ ;
 wire \MuI._1180_ ;
 wire \MuI._1181_ ;
 wire \MuI._1182_ ;
 wire \MuI._1183_ ;
 wire \MuI._1184_ ;
 wire \MuI._1185_ ;
 wire \MuI._1186_ ;
 wire \MuI._1187_ ;
 wire \MuI._1188_ ;
 wire \MuI._1189_ ;
 wire \MuI._1190_ ;
 wire \MuI._1191_ ;
 wire \MuI._1192_ ;
 wire \MuI._1193_ ;
 wire \MuI._1194_ ;
 wire \MuI._1195_ ;
 wire \MuI._1196_ ;
 wire \MuI._1197_ ;
 wire \MuI._1198_ ;
 wire \MuI._1199_ ;
 wire \MuI._1200_ ;
 wire \MuI._1201_ ;
 wire \MuI._1202_ ;
 wire \MuI._1203_ ;
 wire \MuI._1204_ ;
 wire \MuI._1205_ ;
 wire \MuI._1206_ ;
 wire \MuI._1207_ ;
 wire \MuI._1208_ ;
 wire \MuI._1209_ ;
 wire \MuI._1210_ ;
 wire \MuI._1211_ ;
 wire \MuI._1212_ ;
 wire \MuI._1213_ ;
 wire \MuI._1214_ ;
 wire \MuI._1215_ ;
 wire \MuI._1216_ ;
 wire \MuI._1217_ ;
 wire \MuI._1218_ ;
 wire \MuI._1219_ ;
 wire \MuI._1220_ ;
 wire \MuI._1221_ ;
 wire \MuI._1222_ ;
 wire \MuI._1223_ ;
 wire \MuI._1224_ ;
 wire \MuI._1225_ ;
 wire \MuI._1226_ ;
 wire \MuI._1227_ ;
 wire \MuI._1228_ ;
 wire \MuI._1229_ ;
 wire \MuI._1230_ ;
 wire \MuI._1231_ ;
 wire \MuI._1232_ ;
 wire \MuI._1233_ ;
 wire \MuI._1234_ ;
 wire \MuI._1235_ ;
 wire \MuI._1236_ ;
 wire \MuI._1237_ ;
 wire \MuI._1238_ ;
 wire \MuI._1239_ ;
 wire \MuI._1240_ ;
 wire \MuI._1241_ ;
 wire \MuI._1242_ ;
 wire \MuI._1243_ ;
 wire \MuI._1244_ ;
 wire \MuI._1245_ ;
 wire \MuI._1246_ ;
 wire \MuI._1247_ ;
 wire \MuI._1248_ ;
 wire \MuI._1249_ ;
 wire \MuI._1250_ ;
 wire \MuI._1251_ ;
 wire \MuI._1252_ ;
 wire \MuI._1253_ ;
 wire \MuI._1254_ ;
 wire \MuI._1255_ ;
 wire \MuI._1256_ ;
 wire \MuI._1257_ ;
 wire \MuI._1258_ ;
 wire \MuI._1259_ ;
 wire \MuI._1260_ ;
 wire \MuI._1261_ ;
 wire \MuI._1262_ ;
 wire \MuI._1263_ ;
 wire \MuI._1264_ ;
 wire \MuI._1265_ ;
 wire \MuI._1266_ ;
 wire \MuI._1267_ ;
 wire \MuI._1268_ ;
 wire \MuI._1269_ ;
 wire \MuI._1270_ ;
 wire \MuI._1271_ ;
 wire \MuI._1272_ ;
 wire \MuI._1273_ ;
 wire \MuI._1274_ ;
 wire \MuI._1275_ ;
 wire \MuI._1276_ ;
 wire \MuI._1277_ ;
 wire \MuI._1278_ ;
 wire \MuI._1279_ ;
 wire \MuI._1280_ ;
 wire \MuI._1281_ ;
 wire \MuI._1282_ ;
 wire \MuI._1283_ ;
 wire \MuI._1284_ ;
 wire \MuI._1285_ ;
 wire \MuI._1286_ ;
 wire \MuI._1287_ ;
 wire \MuI._1288_ ;
 wire \MuI._1289_ ;
 wire \MuI._1290_ ;
 wire \MuI._1291_ ;
 wire \MuI._1292_ ;
 wire \MuI._1293_ ;
 wire \MuI._1294_ ;
 wire \MuI._1295_ ;
 wire \MuI._1296_ ;
 wire \MuI._1297_ ;
 wire \MuI._1298_ ;
 wire \MuI._1299_ ;
 wire \MuI._1300_ ;
 wire \MuI._1301_ ;
 wire \MuI._1302_ ;
 wire \MuI._1303_ ;
 wire \MuI._1304_ ;
 wire \MuI._1305_ ;
 wire \MuI._1306_ ;
 wire \MuI._1307_ ;
 wire \MuI._1308_ ;
 wire \MuI._1309_ ;
 wire \MuI._1310_ ;
 wire \MuI._1311_ ;
 wire \MuI._1312_ ;
 wire \MuI._1313_ ;
 wire \MuI._1314_ ;
 wire \MuI._1315_ ;
 wire \MuI._1316_ ;
 wire \MuI._1317_ ;
 wire \MuI._1318_ ;
 wire \MuI._1319_ ;
 wire \MuI._1320_ ;
 wire \MuI._1321_ ;
 wire \MuI._1322_ ;
 wire \MuI._1323_ ;
 wire \MuI._1324_ ;
 wire \MuI._1325_ ;
 wire \MuI._1326_ ;
 wire \MuI._1327_ ;
 wire \MuI._1328_ ;
 wire \MuI._1329_ ;
 wire \MuI._1330_ ;
 wire \MuI._1331_ ;
 wire \MuI._1332_ ;
 wire \MuI._1333_ ;
 wire \MuI._1334_ ;
 wire \MuI._1335_ ;
 wire \MuI._1336_ ;
 wire \MuI._1337_ ;
 wire \MuI._1338_ ;
 wire \MuI._1339_ ;
 wire \MuI._1340_ ;
 wire \MuI._1341_ ;
 wire \MuI._1342_ ;
 wire \MuI._1343_ ;
 wire \MuI._1344_ ;
 wire \MuI._1345_ ;
 wire \MuI._1346_ ;
 wire \MuI._1347_ ;
 wire \MuI._1348_ ;
 wire \MuI._1349_ ;
 wire \MuI._1350_ ;
 wire \MuI._1351_ ;
 wire \MuI._1352_ ;
 wire \MuI._1353_ ;
 wire \MuI._1354_ ;
 wire \MuI._1355_ ;
 wire \MuI._1356_ ;
 wire \MuI._1357_ ;
 wire \MuI._1358_ ;
 wire \MuI._1359_ ;
 wire \MuI._1360_ ;
 wire \MuI._1361_ ;
 wire \MuI._1362_ ;
 wire \MuI._1363_ ;
 wire \MuI._1364_ ;
 wire \MuI._1365_ ;
 wire \MuI._1366_ ;
 wire \MuI._1367_ ;
 wire \MuI._1368_ ;
 wire \MuI._1369_ ;
 wire \MuI._1370_ ;
 wire \MuI._1371_ ;
 wire \MuI._1372_ ;
 wire \MuI._1373_ ;
 wire \MuI._1374_ ;
 wire \MuI._1375_ ;
 wire \MuI._1376_ ;
 wire \MuI._1377_ ;
 wire \MuI._1378_ ;
 wire \MuI._1379_ ;
 wire \MuI._1380_ ;
 wire \MuI._1381_ ;
 wire \MuI._1382_ ;
 wire \MuI._1383_ ;
 wire \MuI._1384_ ;
 wire \MuI._1385_ ;
 wire \MuI._1386_ ;
 wire \MuI._1387_ ;
 wire \MuI._1388_ ;
 wire \MuI._1389_ ;
 wire \MuI._1390_ ;
 wire \MuI._1391_ ;
 wire \MuI._1392_ ;
 wire \MuI._1393_ ;
 wire \MuI._1394_ ;
 wire \MuI._1395_ ;
 wire \MuI._1396_ ;
 wire \MuI._1397_ ;
 wire \MuI._1398_ ;
 wire \MuI._1399_ ;
 wire \MuI._1400_ ;
 wire \MuI._1401_ ;
 wire \MuI._1402_ ;
 wire \MuI._1403_ ;
 wire \MuI._1404_ ;
 wire \MuI._1405_ ;
 wire \MuI._1406_ ;
 wire \MuI._1407_ ;
 wire \MuI._1408_ ;
 wire \MuI._1409_ ;
 wire \MuI._1410_ ;
 wire \MuI._1411_ ;
 wire \MuI._1412_ ;
 wire \MuI._1413_ ;
 wire \MuI._1414_ ;
 wire \MuI._1415_ ;
 wire \MuI._1416_ ;
 wire \MuI._1417_ ;
 wire \MuI._1418_ ;
 wire \MuI._1419_ ;
 wire \MuI._1420_ ;
 wire \MuI._1421_ ;
 wire \MuI._1422_ ;
 wire \MuI._1423_ ;
 wire \MuI._1424_ ;
 wire \MuI._1425_ ;
 wire \MuI._1426_ ;
 wire \MuI._1427_ ;
 wire \MuI._1428_ ;
 wire \MuI._1429_ ;
 wire \MuI._1430_ ;
 wire \MuI._1431_ ;
 wire \MuI._1432_ ;
 wire \MuI._1433_ ;
 wire \MuI._1434_ ;
 wire \MuI._1435_ ;
 wire \MuI._1436_ ;
 wire \MuI._1437_ ;
 wire \MuI._1438_ ;
 wire \MuI._1439_ ;
 wire \MuI._1440_ ;
 wire \MuI._1441_ ;
 wire \MuI._1442_ ;
 wire \MuI._1443_ ;
 wire \MuI._1444_ ;
 wire \MuI._1445_ ;
 wire \MuI._1446_ ;
 wire \MuI._1447_ ;
 wire \MuI._1448_ ;
 wire \MuI._1449_ ;
 wire \MuI._1450_ ;
 wire \MuI._1451_ ;
 wire \MuI._1452_ ;
 wire \MuI._1453_ ;
 wire \MuI._1454_ ;
 wire \MuI._1455_ ;
 wire \MuI._1456_ ;
 wire \MuI._1457_ ;
 wire \MuI._1458_ ;
 wire \MuI._1459_ ;
 wire \MuI._1460_ ;
 wire \MuI._1461_ ;
 wire \MuI._1462_ ;
 wire \MuI._1463_ ;
 wire \MuI._1464_ ;
 wire \MuI._1465_ ;
 wire \MuI._1466_ ;
 wire \MuI._1467_ ;
 wire \MuI._1468_ ;
 wire \MuI._1469_ ;
 wire \MuI._1470_ ;
 wire \MuI._1471_ ;
 wire \MuI._1472_ ;
 wire \MuI._1473_ ;
 wire \MuI._1474_ ;
 wire \MuI._1475_ ;
 wire \MuI._1476_ ;
 wire \MuI._1477_ ;
 wire \MuI._1478_ ;
 wire \MuI._1479_ ;
 wire \MuI._1480_ ;
 wire \MuI._1481_ ;
 wire \MuI._1482_ ;
 wire \MuI._1483_ ;
 wire \MuI._1484_ ;
 wire \MuI._1485_ ;
 wire \MuI._1486_ ;
 wire \MuI._1487_ ;
 wire \MuI._1488_ ;
 wire \MuI._1489_ ;
 wire \MuI._1490_ ;
 wire \MuI._1491_ ;
 wire \MuI._1492_ ;
 wire \MuI._1493_ ;
 wire \MuI._1494_ ;
 wire \MuI._1495_ ;
 wire \MuI._1496_ ;
 wire \MuI._1497_ ;
 wire \MuI._1498_ ;
 wire \MuI._1499_ ;
 wire \MuI._1500_ ;
 wire \MuI._1501_ ;
 wire \MuI._1502_ ;
 wire \MuI._1503_ ;
 wire \MuI._1504_ ;
 wire \MuI._1505_ ;
 wire \MuI._1506_ ;
 wire \MuI._1507_ ;
 wire \MuI._1508_ ;
 wire \MuI._1509_ ;
 wire \MuI._1510_ ;
 wire \MuI._1511_ ;
 wire \MuI._1512_ ;
 wire \MuI._1513_ ;
 wire \MuI._1514_ ;
 wire \MuI._1515_ ;
 wire \MuI._1516_ ;
 wire \MuI._1517_ ;
 wire \MuI._1518_ ;
 wire \MuI._1519_ ;
 wire \MuI._1520_ ;
 wire \MuI._1521_ ;
 wire \MuI._1522_ ;
 wire \MuI._1523_ ;
 wire \MuI._1524_ ;
 wire \MuI._1525_ ;
 wire \MuI._1526_ ;
 wire \MuI._1527_ ;
 wire \MuI._1528_ ;
 wire \MuI._1529_ ;
 wire \MuI._1530_ ;
 wire \MuI._1531_ ;
 wire \MuI._1532_ ;
 wire \MuI._1533_ ;
 wire \MuI._1534_ ;
 wire \MuI._1535_ ;
 wire \MuI._1536_ ;
 wire \MuI._1537_ ;
 wire \MuI._1538_ ;
 wire \MuI._1539_ ;
 wire \MuI._1540_ ;
 wire \MuI._1541_ ;
 wire \MuI._1542_ ;
 wire \MuI._1543_ ;
 wire \MuI._1544_ ;
 wire \MuI._1545_ ;
 wire \MuI._1546_ ;
 wire \MuI._1547_ ;
 wire \MuI._1548_ ;
 wire \MuI._1549_ ;
 wire \MuI._1550_ ;
 wire \MuI._1551_ ;
 wire \MuI._1552_ ;
 wire \MuI._1553_ ;
 wire \MuI._1554_ ;
 wire \MuI._1555_ ;
 wire \MuI._1556_ ;
 wire \MuI._1557_ ;
 wire \MuI._1558_ ;
 wire \MuI._1559_ ;
 wire \MuI._1560_ ;
 wire \MuI._1561_ ;
 wire \MuI._1562_ ;
 wire \MuI._1563_ ;
 wire \MuI._1564_ ;
 wire \MuI._1565_ ;
 wire \MuI._1566_ ;
 wire \MuI._1567_ ;
 wire \MuI._1568_ ;
 wire \MuI._1569_ ;
 wire \MuI._1570_ ;
 wire \MuI._1571_ ;
 wire \MuI._1572_ ;
 wire \MuI._1573_ ;
 wire \MuI._1574_ ;
 wire \MuI._1575_ ;
 wire \MuI._1576_ ;
 wire \MuI._1577_ ;
 wire \MuI._1578_ ;
 wire \MuI._1579_ ;
 wire \MuI._1580_ ;
 wire \MuI._1581_ ;
 wire \MuI._1582_ ;
 wire \MuI._1583_ ;
 wire \MuI._1584_ ;
 wire \MuI._1585_ ;
 wire \MuI._1586_ ;
 wire \MuI._1587_ ;
 wire \MuI._1588_ ;
 wire \MuI._1589_ ;
 wire \MuI._1590_ ;
 wire \MuI._1591_ ;
 wire \MuI._1592_ ;
 wire \MuI._1593_ ;
 wire \MuI._1594_ ;
 wire \MuI._1595_ ;
 wire \MuI._1596_ ;
 wire \MuI._1597_ ;
 wire \MuI._1598_ ;
 wire \MuI._1599_ ;
 wire \MuI._1600_ ;
 wire \MuI._1601_ ;
 wire \MuI._1602_ ;
 wire \MuI._1603_ ;
 wire \MuI._1604_ ;
 wire \MuI._1605_ ;
 wire \MuI._1606_ ;
 wire \MuI._1607_ ;
 wire \MuI._1608_ ;
 wire \MuI._1609_ ;
 wire \MuI._1610_ ;
 wire \MuI._1611_ ;
 wire \MuI._1612_ ;
 wire \MuI._1613_ ;
 wire \MuI._1614_ ;
 wire \MuI._1615_ ;
 wire \MuI._1616_ ;
 wire \MuI._1617_ ;
 wire \MuI._1618_ ;
 wire \MuI._1619_ ;
 wire \MuI._1620_ ;
 wire \MuI._1621_ ;
 wire \MuI._1622_ ;
 wire \MuI._1623_ ;
 wire \MuI._1624_ ;
 wire \MuI._1625_ ;
 wire \MuI._1626_ ;
 wire \MuI._1627_ ;
 wire \MuI._1628_ ;
 wire \MuI._1629_ ;
 wire \MuI._1630_ ;
 wire \MuI._1631_ ;
 wire \MuI._1632_ ;
 wire \MuI._1633_ ;
 wire \MuI._1634_ ;
 wire \MuI._1635_ ;
 wire \MuI._1636_ ;
 wire \MuI._1637_ ;
 wire \MuI._1638_ ;
 wire \MuI._1639_ ;
 wire \MuI._1640_ ;
 wire \MuI._1641_ ;
 wire \MuI._1642_ ;
 wire \MuI._1643_ ;
 wire \MuI._1644_ ;
 wire \MuI._1645_ ;
 wire \MuI._1646_ ;
 wire \MuI._1647_ ;
 wire \MuI._1648_ ;
 wire \MuI._1649_ ;
 wire \MuI._1650_ ;
 wire \MuI._1651_ ;
 wire \MuI._1652_ ;
 wire \MuI._1653_ ;
 wire \MuI._1654_ ;
 wire \MuI._1655_ ;
 wire \MuI._1656_ ;
 wire \MuI._1657_ ;
 wire \MuI._1658_ ;
 wire \MuI._1659_ ;
 wire \MuI._1660_ ;
 wire \MuI._1661_ ;
 wire \MuI._1662_ ;
 wire \MuI._1663_ ;
 wire \MuI._1664_ ;
 wire \MuI._1665_ ;
 wire \MuI._1666_ ;
 wire \MuI._1667_ ;
 wire \MuI._1668_ ;
 wire \MuI._1669_ ;
 wire \MuI._1670_ ;
 wire \MuI._1671_ ;
 wire \MuI._1672_ ;
 wire \MuI._1673_ ;
 wire \MuI._1674_ ;
 wire \MuI._1675_ ;
 wire \MuI._1676_ ;
 wire \MuI._1677_ ;
 wire \MuI._1678_ ;
 wire \MuI._1679_ ;
 wire \MuI._1680_ ;
 wire \MuI._1681_ ;
 wire \MuI._1682_ ;
 wire \MuI._1683_ ;
 wire \MuI._1684_ ;
 wire \MuI._1685_ ;
 wire \MuI._1686_ ;
 wire \MuI._1687_ ;
 wire \MuI._1688_ ;
 wire \MuI._1689_ ;
 wire \MuI._1690_ ;
 wire \MuI._1691_ ;
 wire \MuI._1692_ ;
 wire \MuI._1693_ ;
 wire \MuI._1694_ ;
 wire \MuI._1695_ ;
 wire \MuI._1696_ ;
 wire \MuI._1697_ ;
 wire \MuI._1698_ ;
 wire \MuI._1699_ ;
 wire \MuI._1700_ ;
 wire \MuI._1701_ ;
 wire \MuI._1702_ ;
 wire \MuI._1703_ ;
 wire \MuI._1704_ ;
 wire \MuI._1705_ ;
 wire \MuI._1706_ ;
 wire \MuI._1707_ ;
 wire \MuI._1708_ ;
 wire \MuI._1709_ ;
 wire \MuI._1710_ ;
 wire \MuI._1711_ ;
 wire \MuI._1712_ ;
 wire \MuI._1713_ ;
 wire \MuI._1714_ ;
 wire \MuI._1715_ ;
 wire \MuI._1716_ ;
 wire \MuI._1717_ ;
 wire \MuI._1718_ ;
 wire \MuI._1719_ ;
 wire \MuI._1720_ ;
 wire \MuI._1721_ ;
 wire \MuI._1722_ ;
 wire \MuI._1723_ ;
 wire \MuI._1724_ ;
 wire \MuI._1725_ ;
 wire \MuI._1726_ ;
 wire \MuI._1727_ ;
 wire \MuI._1728_ ;
 wire \MuI._1729_ ;
 wire \MuI._1730_ ;
 wire \MuI._1731_ ;
 wire \MuI._1732_ ;
 wire \MuI._1733_ ;
 wire \MuI._1734_ ;
 wire \MuI._1735_ ;
 wire \MuI._1736_ ;
 wire \MuI._1737_ ;
 wire \MuI._1738_ ;
 wire \MuI._1739_ ;
 wire \MuI._1740_ ;
 wire \MuI._1741_ ;
 wire \MuI._1742_ ;
 wire \MuI._1743_ ;
 wire \MuI._1744_ ;
 wire \MuI._1745_ ;
 wire \MuI._1746_ ;
 wire \MuI._1747_ ;
 wire \MuI._1748_ ;
 wire \MuI._1749_ ;
 wire \MuI._1750_ ;
 wire \MuI._1751_ ;
 wire \MuI._1752_ ;
 wire \MuI._1753_ ;
 wire \MuI._1754_ ;
 wire \MuI._1755_ ;
 wire \MuI._1756_ ;
 wire \MuI._1757_ ;
 wire \MuI._1758_ ;
 wire \MuI._1759_ ;
 wire \MuI._1760_ ;
 wire \MuI._1761_ ;
 wire \MuI._1762_ ;
 wire \MuI._1763_ ;
 wire \MuI._1764_ ;
 wire \MuI._1765_ ;
 wire \MuI._1766_ ;
 wire \MuI._1767_ ;
 wire \MuI._1768_ ;
 wire \MuI._1769_ ;
 wire \MuI._1770_ ;
 wire \MuI._1771_ ;
 wire \MuI._1772_ ;
 wire \MuI._1773_ ;
 wire \MuI._1774_ ;
 wire \MuI._1775_ ;
 wire \MuI._1776_ ;
 wire \MuI._1777_ ;
 wire \MuI._1778_ ;
 wire \MuI._1779_ ;
 wire \MuI._1780_ ;
 wire \MuI._1781_ ;
 wire \MuI._1782_ ;
 wire \MuI._1783_ ;
 wire \MuI._1784_ ;
 wire \MuI._1785_ ;
 wire \MuI._1786_ ;
 wire \MuI._1787_ ;
 wire \MuI._1788_ ;
 wire \MuI._1789_ ;
 wire \MuI._1790_ ;
 wire \MuI._1791_ ;
 wire \MuI._1792_ ;
 wire \MuI._1793_ ;
 wire \MuI._1794_ ;
 wire \MuI._1795_ ;
 wire \MuI._1796_ ;
 wire \MuI._1797_ ;
 wire \MuI._1798_ ;
 wire \MuI._1799_ ;
 wire \MuI._1800_ ;
 wire \MuI._1801_ ;
 wire \MuI._1802_ ;
 wire \MuI._1803_ ;
 wire \MuI._1804_ ;
 wire \MuI._1805_ ;
 wire \MuI._1806_ ;
 wire \MuI._1807_ ;
 wire \MuI._1808_ ;
 wire \MuI._1809_ ;
 wire \MuI._1810_ ;
 wire \MuI._1811_ ;
 wire \MuI._1812_ ;
 wire \MuI._1813_ ;
 wire \MuI._1814_ ;
 wire \MuI._1815_ ;
 wire \MuI._1816_ ;
 wire \MuI._1817_ ;
 wire \MuI._1818_ ;
 wire \MuI._1819_ ;
 wire \MuI._1820_ ;
 wire \MuI._1821_ ;
 wire \MuI._1822_ ;
 wire \MuI._1823_ ;
 wire \MuI._1824_ ;
 wire \MuI._1825_ ;
 wire \MuI._1826_ ;
 wire \MuI._1827_ ;
 wire \MuI._1828_ ;
 wire \MuI._1829_ ;
 wire \MuI._1830_ ;
 wire \MuI._1831_ ;
 wire \MuI._1832_ ;
 wire \MuI._1833_ ;
 wire \MuI._1834_ ;
 wire \MuI._1835_ ;
 wire \MuI._1836_ ;
 wire \MuI._1837_ ;
 wire \MuI._1838_ ;
 wire \MuI._1839_ ;
 wire \MuI._1840_ ;
 wire \MuI._1841_ ;
 wire \MuI._1842_ ;
 wire \MuI._1843_ ;
 wire \MuI._1844_ ;
 wire \MuI._1845_ ;
 wire \MuI._1846_ ;
 wire \MuI._1847_ ;
 wire \MuI._1848_ ;
 wire \MuI._1849_ ;
 wire \MuI._1850_ ;
 wire \MuI._1851_ ;
 wire \MuI._1852_ ;
 wire \MuI._1853_ ;
 wire \MuI._1854_ ;
 wire \MuI._1855_ ;
 wire \MuI._1856_ ;
 wire \MuI._1857_ ;
 wire \MuI._1858_ ;
 wire \MuI._1859_ ;
 wire \MuI._1860_ ;
 wire \MuI._1861_ ;
 wire \MuI._1862_ ;
 wire \MuI._1863_ ;
 wire \MuI._1864_ ;
 wire \MuI._1865_ ;
 wire \MuI._1866_ ;
 wire \MuI._1867_ ;
 wire \MuI._1868_ ;
 wire \MuI._1869_ ;
 wire \MuI._1870_ ;
 wire \MuI._1871_ ;
 wire \MuI._1872_ ;
 wire \MuI._1873_ ;
 wire \MuI._1874_ ;
 wire \MuI._1875_ ;
 wire \MuI._1876_ ;
 wire \MuI._1877_ ;
 wire \MuI._1878_ ;
 wire \MuI._1879_ ;
 wire \MuI._1880_ ;
 wire \MuI._1881_ ;
 wire \MuI._1882_ ;
 wire \MuI._1883_ ;
 wire \MuI._1884_ ;
 wire \MuI._1885_ ;
 wire \MuI._1886_ ;
 wire \MuI._1887_ ;
 wire \MuI._1888_ ;
 wire \MuI._1889_ ;
 wire \MuI._1890_ ;
 wire \MuI._1891_ ;
 wire \MuI._1892_ ;
 wire \MuI._1893_ ;
 wire \MuI._1894_ ;
 wire \MuI._1895_ ;
 wire \MuI._1896_ ;
 wire \MuI._1897_ ;
 wire \MuI._1898_ ;
 wire \MuI._1899_ ;
 wire \MuI._1900_ ;
 wire \MuI._1901_ ;
 wire \MuI._1902_ ;
 wire \MuI._1903_ ;
 wire \MuI._1904_ ;
 wire \MuI._1905_ ;
 wire \MuI._1906_ ;
 wire \MuI._1907_ ;
 wire \MuI._1908_ ;
 wire \MuI._1909_ ;
 wire \MuI._1910_ ;
 wire \MuI._1911_ ;
 wire \MuI._1912_ ;
 wire \MuI._1913_ ;
 wire \MuI._1914_ ;
 wire \MuI._1915_ ;
 wire \MuI._1916_ ;
 wire \MuI._1917_ ;
 wire \MuI._1918_ ;
 wire \MuI._1919_ ;
 wire \MuI._1920_ ;
 wire \MuI._1921_ ;
 wire \MuI._1922_ ;
 wire \MuI._1923_ ;
 wire \MuI._1924_ ;
 wire \MuI._1925_ ;
 wire \MuI._1926_ ;
 wire \MuI._1927_ ;
 wire \MuI._1928_ ;
 wire \MuI._1929_ ;
 wire \MuI._1930_ ;
 wire \MuI._1931_ ;
 wire \MuI._1932_ ;
 wire \MuI._1933_ ;
 wire \MuI._1934_ ;
 wire \MuI._1935_ ;
 wire \MuI._1936_ ;
 wire \MuI._1937_ ;
 wire \MuI._1938_ ;
 wire \MuI._1939_ ;
 wire \MuI._1940_ ;
 wire \MuI._1941_ ;
 wire \MuI._1942_ ;
 wire \MuI._1943_ ;
 wire \MuI._1944_ ;
 wire \MuI._1945_ ;
 wire \MuI._1946_ ;
 wire \MuI._1947_ ;
 wire \MuI._1948_ ;
 wire \MuI._1949_ ;
 wire \MuI._1950_ ;
 wire \MuI._1951_ ;
 wire \MuI._1952_ ;
 wire \MuI._1953_ ;
 wire \MuI._1954_ ;
 wire \MuI._1955_ ;
 wire \MuI._1956_ ;
 wire \MuI._1957_ ;
 wire \MuI._1958_ ;
 wire \MuI._1959_ ;
 wire \MuI._1960_ ;
 wire \MuI._1961_ ;
 wire \MuI._1962_ ;
 wire \MuI._1963_ ;
 wire \MuI._1964_ ;
 wire \MuI._1965_ ;
 wire \MuI._1966_ ;
 wire \MuI._1967_ ;
 wire \MuI._1968_ ;
 wire \MuI._1969_ ;
 wire \MuI._1970_ ;
 wire \MuI._1971_ ;
 wire \MuI._1972_ ;
 wire \MuI._1973_ ;
 wire \MuI._1974_ ;
 wire \MuI._1975_ ;
 wire \MuI._1976_ ;
 wire \MuI._1977_ ;
 wire \MuI._1978_ ;
 wire \MuI._1979_ ;
 wire \MuI._1980_ ;
 wire \MuI._1981_ ;
 wire \MuI._1982_ ;
 wire \MuI._1983_ ;
 wire \MuI._1984_ ;
 wire \MuI._1985_ ;
 wire \MuI._1986_ ;
 wire \MuI._1987_ ;
 wire \MuI._1988_ ;
 wire \MuI._1989_ ;
 wire \MuI._1990_ ;
 wire \MuI._1991_ ;
 wire \MuI._1992_ ;
 wire \MuI._1993_ ;
 wire \MuI._1994_ ;
 wire \MuI._1995_ ;
 wire \MuI._1996_ ;
 wire \MuI._1997_ ;
 wire \MuI._1998_ ;
 wire \MuI._1999_ ;
 wire \MuI._2000_ ;
 wire \MuI._2001_ ;
 wire \MuI._2002_ ;
 wire \MuI._2003_ ;
 wire \MuI._2004_ ;
 wire \MuI._2005_ ;
 wire \MuI._2006_ ;
 wire \MuI._2007_ ;
 wire \MuI._2008_ ;
 wire \MuI._2009_ ;
 wire \MuI._2010_ ;
 wire \MuI._2011_ ;
 wire \MuI._2012_ ;
 wire \MuI._2013_ ;
 wire \MuI._2014_ ;
 wire \MuI._2015_ ;
 wire \MuI._2016_ ;
 wire \MuI._2017_ ;
 wire \MuI._2018_ ;
 wire \MuI._2019_ ;
 wire \MuI._2020_ ;
 wire \MuI._2021_ ;
 wire \MuI._2022_ ;
 wire \MuI._2023_ ;
 wire \MuI._2024_ ;
 wire \MuI._2025_ ;
 wire \MuI._2026_ ;
 wire \MuI._2027_ ;
 wire \MuI._2028_ ;
 wire \MuI._2029_ ;
 wire \MuI._2030_ ;
 wire \MuI._2031_ ;
 wire \MuI._2032_ ;
 wire \MuI._2033_ ;
 wire \MuI._2034_ ;
 wire \MuI._2035_ ;
 wire \MuI._2036_ ;
 wire \MuI._2037_ ;
 wire \MuI._2038_ ;
 wire \MuI._2039_ ;
 wire \MuI._2040_ ;
 wire \MuI._2041_ ;
 wire \MuI._2042_ ;
 wire \MuI._2043_ ;
 wire \MuI._2044_ ;
 wire \MuI._2045_ ;
 wire \MuI._2046_ ;
 wire \MuI._2047_ ;
 wire \MuI._2048_ ;
 wire \MuI._2049_ ;
 wire \MuI._2050_ ;
 wire \MuI._2051_ ;
 wire \MuI._2052_ ;
 wire \MuI._2053_ ;
 wire \MuI._2054_ ;
 wire \MuI._2055_ ;
 wire \MuI._2056_ ;
 wire \MuI._2057_ ;
 wire \MuI._2058_ ;
 wire \MuI._2059_ ;
 wire \MuI._2060_ ;
 wire \MuI._2061_ ;
 wire \MuI._2062_ ;
 wire \MuI._2063_ ;
 wire \MuI._2064_ ;
 wire \MuI._2065_ ;
 wire \MuI._2066_ ;
 wire \MuI._2067_ ;
 wire \MuI._2068_ ;
 wire \MuI._2069_ ;
 wire \MuI._2070_ ;
 wire \MuI._2071_ ;
 wire \MuI._2072_ ;
 wire \MuI._2073_ ;
 wire \MuI._2074_ ;
 wire \MuI._2075_ ;
 wire \MuI._2076_ ;
 wire \MuI._2077_ ;
 wire \MuI._2078_ ;
 wire \MuI._2079_ ;
 wire \MuI._2080_ ;
 wire \MuI._2081_ ;
 wire \MuI._2082_ ;
 wire \MuI._2083_ ;
 wire \MuI._2084_ ;
 wire \MuI._2085_ ;
 wire \MuI._2086_ ;
 wire \MuI._2087_ ;
 wire \MuI._2088_ ;
 wire \MuI._2089_ ;
 wire \MuI._2090_ ;
 wire \MuI._2091_ ;
 wire \MuI._2092_ ;
 wire \MuI._2093_ ;
 wire \MuI._2094_ ;
 wire \MuI._2095_ ;
 wire \MuI._2096_ ;
 wire \MuI._2097_ ;
 wire \MuI._2098_ ;
 wire \MuI._2099_ ;
 wire \MuI._2100_ ;
 wire \MuI._2101_ ;
 wire \MuI._2102_ ;
 wire \MuI._2103_ ;
 wire \MuI._2104_ ;
 wire \MuI._2105_ ;
 wire \MuI._2106_ ;
 wire \MuI._2107_ ;
 wire \MuI._2108_ ;
 wire \MuI._2109_ ;
 wire \MuI._2110_ ;
 wire \MuI._2111_ ;
 wire \MuI._2112_ ;
 wire \MuI._2113_ ;
 wire \MuI._2114_ ;
 wire \MuI._2115_ ;
 wire \MuI._2116_ ;
 wire \MuI._2117_ ;
 wire \MuI._2118_ ;
 wire \MuI._2119_ ;
 wire \MuI._2120_ ;
 wire \MuI._2121_ ;
 wire \MuI._2122_ ;
 wire \MuI._2123_ ;
 wire \MuI._2124_ ;
 wire \MuI._2125_ ;
 wire \MuI._2126_ ;
 wire \MuI._2127_ ;
 wire \MuI._2128_ ;
 wire \MuI._2129_ ;
 wire \MuI._2130_ ;
 wire \MuI._2131_ ;
 wire \MuI._2132_ ;
 wire \MuI._2133_ ;
 wire \MuI._2134_ ;
 wire \MuI._2135_ ;
 wire \MuI._2136_ ;
 wire \MuI._2137_ ;
 wire \MuI._2138_ ;
 wire \MuI._2139_ ;
 wire \MuI._2140_ ;
 wire \MuI._2141_ ;
 wire \MuI._2142_ ;
 wire \MuI._2143_ ;
 wire \MuI._2144_ ;
 wire \MuI._2145_ ;
 wire \MuI._2146_ ;
 wire \MuI._2147_ ;
 wire \MuI._2148_ ;
 wire \MuI._2149_ ;
 wire \MuI._2150_ ;
 wire \MuI._2151_ ;
 wire \MuI._2152_ ;
 wire \MuI._2153_ ;
 wire \MuI._2154_ ;
 wire \MuI._2155_ ;
 wire \MuI._2156_ ;
 wire \MuI._2157_ ;
 wire \MuI._2158_ ;
 wire \MuI._2159_ ;
 wire \MuI._2160_ ;
 wire \MuI._2161_ ;
 wire \MuI._2162_ ;
 wire \MuI._2163_ ;
 wire \MuI._2164_ ;
 wire \MuI._2165_ ;
 wire \MuI._2166_ ;
 wire \MuI._2167_ ;
 wire \MuI._2168_ ;
 wire \MuI._2169_ ;
 wire \MuI._2170_ ;
 wire \MuI._2171_ ;
 wire \MuI._2172_ ;
 wire \MuI._2173_ ;
 wire \MuI._2174_ ;
 wire \MuI._2175_ ;
 wire \MuI._2176_ ;
 wire \MuI._2177_ ;
 wire \MuI._2178_ ;
 wire \MuI._2179_ ;
 wire \MuI._2180_ ;
 wire \MuI._2181_ ;
 wire \MuI._2182_ ;
 wire \MuI._2183_ ;
 wire \MuI._2184_ ;
 wire \MuI._2185_ ;
 wire \MuI._2186_ ;
 wire \MuI._2187_ ;
 wire \MuI._2188_ ;
 wire \MuI._2189_ ;
 wire \MuI._2190_ ;
 wire \MuI._2191_ ;
 wire \MuI._2192_ ;
 wire \MuI._2193_ ;
 wire \MuI._2194_ ;
 wire \MuI._2195_ ;
 wire \MuI._2196_ ;
 wire \MuI._2197_ ;
 wire \MuI._2198_ ;
 wire \MuI._2199_ ;
 wire \MuI._2200_ ;
 wire \MuI._2201_ ;
 wire \MuI._2202_ ;
 wire \MuI._2203_ ;
 wire \MuI._2204_ ;
 wire \MuI._2205_ ;
 wire \MuI._2206_ ;
 wire \MuI._2207_ ;
 wire \MuI._2208_ ;
 wire \MuI._2209_ ;
 wire \MuI._2210_ ;
 wire \MuI._2211_ ;
 wire \MuI._2212_ ;
 wire \MuI._2213_ ;
 wire \MuI._2214_ ;
 wire \MuI._2215_ ;
 wire \MuI._2216_ ;
 wire \MuI._2217_ ;
 wire \MuI._2218_ ;
 wire \MuI._2219_ ;
 wire \MuI._2220_ ;
 wire \MuI._2221_ ;
 wire \MuI._2222_ ;
 wire \MuI._2223_ ;
 wire \MuI._2224_ ;
 wire \MuI._2225_ ;
 wire \MuI._2226_ ;
 wire \MuI._2227_ ;
 wire \MuI._2228_ ;
 wire \MuI._2229_ ;
 wire \MuI._2230_ ;
 wire \MuI._2231_ ;
 wire \MuI._2232_ ;
 wire \MuI._2233_ ;
 wire \MuI._2234_ ;
 wire \MuI._2235_ ;
 wire \MuI._2236_ ;
 wire \MuI._2237_ ;
 wire \MuI._2238_ ;
 wire \MuI._2239_ ;
 wire \MuI._2240_ ;
 wire \MuI._2241_ ;
 wire \MuI._2242_ ;
 wire \MuI._2243_ ;
 wire \MuI._2244_ ;
 wire \MuI._2245_ ;
 wire \MuI._2246_ ;
 wire \MuI._2247_ ;
 wire \MuI._2248_ ;
 wire \MuI._2249_ ;
 wire \MuI._2250_ ;
 wire \MuI._2251_ ;
 wire \MuI._2252_ ;
 wire \MuI._2253_ ;
 wire \MuI._2254_ ;
 wire \MuI._2255_ ;
 wire \MuI._2256_ ;
 wire \MuI._2257_ ;
 wire \MuI._2258_ ;
 wire \MuI._2259_ ;
 wire \MuI._2260_ ;
 wire \MuI._2261_ ;
 wire \MuI._2262_ ;
 wire \MuI._2263_ ;
 wire \MuI._2264_ ;
 wire \MuI._2265_ ;
 wire \MuI._2266_ ;
 wire \MuI._2267_ ;
 wire \MuI._2268_ ;
 wire \MuI._2269_ ;
 wire \MuI._2270_ ;
 wire \MuI._2271_ ;
 wire \MuI._2272_ ;
 wire \MuI._2273_ ;
 wire \MuI._2274_ ;
 wire \MuI._2275_ ;
 wire \MuI._2276_ ;
 wire \MuI._2277_ ;
 wire \MuI._2278_ ;
 wire \MuI._2279_ ;
 wire \MuI._2280_ ;
 wire \MuI._2281_ ;
 wire \MuI._2282_ ;
 wire \MuI._2283_ ;
 wire \MuI._2284_ ;
 wire \MuI._2285_ ;
 wire \MuI._2286_ ;
 wire \MuI._2287_ ;
 wire \MuI._2288_ ;
 wire \MuI._2289_ ;
 wire \MuI._2290_ ;
 wire \MuI._2291_ ;
 wire \MuI._2292_ ;
 wire \MuI._2293_ ;
 wire \MuI._2294_ ;
 wire \MuI._2295_ ;
 wire \MuI._2296_ ;
 wire \MuI._2297_ ;
 wire \MuI._2298_ ;
 wire \MuI._2299_ ;
 wire \MuI._2300_ ;
 wire \MuI._2301_ ;
 wire \MuI._2302_ ;
 wire \MuI._2303_ ;
 wire \MuI._2304_ ;
 wire \MuI._2305_ ;
 wire \MuI._2306_ ;
 wire \MuI._2307_ ;
 wire \MuI._2308_ ;
 wire \MuI._2309_ ;
 wire \MuI._2310_ ;
 wire \MuI._2311_ ;
 wire \MuI._2312_ ;
 wire \MuI._2313_ ;
 wire \MuI._2314_ ;
 wire \MuI._2315_ ;
 wire \MuI._2316_ ;
 wire \MuI._2317_ ;
 wire \MuI._2318_ ;
 wire \MuI._2319_ ;
 wire \MuI._2320_ ;
 wire \MuI._2321_ ;
 wire \MuI._2322_ ;
 wire \MuI._2323_ ;
 wire \MuI._2324_ ;
 wire \MuI._2325_ ;
 wire \MuI._2326_ ;
 wire \MuI._2327_ ;
 wire \MuI._2328_ ;
 wire \MuI._2329_ ;
 wire \MuI._2330_ ;
 wire \MuI._2331_ ;
 wire \MuI._2332_ ;
 wire \MuI._2333_ ;
 wire \MuI._2334_ ;
 wire \MuI._2335_ ;
 wire \MuI._2336_ ;
 wire \MuI._2337_ ;
 wire \MuI._2338_ ;
 wire \MuI._2339_ ;
 wire \MuI._2340_ ;
 wire \MuI._2341_ ;
 wire \MuI._2342_ ;
 wire \MuI._2343_ ;
 wire \MuI._2344_ ;
 wire \MuI._2345_ ;
 wire \MuI._2346_ ;
 wire \MuI._2347_ ;
 wire \MuI._2348_ ;
 wire \MuI._2349_ ;
 wire \MuI._2350_ ;
 wire \MuI._2351_ ;
 wire \MuI._2352_ ;
 wire \MuI._2353_ ;
 wire \MuI._2354_ ;
 wire \MuI._2355_ ;
 wire \MuI._2356_ ;
 wire \MuI._2357_ ;
 wire \MuI._2358_ ;
 wire \MuI._2359_ ;
 wire \MuI._2360_ ;
 wire \MuI._2361_ ;
 wire \MuI._2362_ ;
 wire \MuI._2363_ ;
 wire \MuI._2364_ ;
 wire \MuI._2365_ ;
 wire \MuI._2366_ ;
 wire \MuI._2367_ ;
 wire \MuI._2368_ ;
 wire \MuI._2369_ ;
 wire \MuI._2370_ ;
 wire \MuI._2371_ ;
 wire \MuI._2372_ ;
 wire \MuI._2373_ ;
 wire \MuI._2374_ ;
 wire \MuI._2375_ ;
 wire \MuI._2376_ ;
 wire \MuI._2377_ ;
 wire \MuI._2378_ ;
 wire \MuI._2379_ ;
 wire \MuI._2380_ ;
 wire \MuI._2381_ ;
 wire \MuI._2382_ ;
 wire \MuI._2383_ ;
 wire \MuI._2384_ ;
 wire \MuI._2385_ ;
 wire \MuI._2386_ ;
 wire \MuI._2387_ ;
 wire \MuI._2388_ ;
 wire \MuI._2389_ ;
 wire \MuI._2390_ ;
 wire \MuI._2391_ ;
 wire \MuI._2392_ ;
 wire \MuI._2393_ ;
 wire \MuI._2394_ ;
 wire \MuI._2395_ ;
 wire \MuI._2396_ ;
 wire \MuI._2397_ ;
 wire \MuI._2398_ ;
 wire \MuI._2399_ ;
 wire \MuI._2400_ ;
 wire \MuI._2401_ ;
 wire \MuI._2402_ ;
 wire \MuI._2403_ ;
 wire \MuI._2404_ ;
 wire \MuI._2405_ ;
 wire \MuI._2406_ ;
 wire \MuI._2407_ ;
 wire \MuI._2408_ ;
 wire \MuI._2409_ ;
 wire \MuI._2410_ ;
 wire \MuI._2411_ ;
 wire \MuI._2412_ ;
 wire \MuI._2413_ ;
 wire \MuI._2414_ ;
 wire \MuI._2415_ ;
 wire \MuI._2416_ ;
 wire \MuI._2417_ ;
 wire \MuI._2418_ ;
 wire \MuI._2419_ ;
 wire \MuI._2420_ ;
 wire \MuI._2421_ ;
 wire \MuI._2422_ ;
 wire \MuI._2423_ ;
 wire \MuI._2424_ ;
 wire \MuI._2425_ ;
 wire \MuI._2426_ ;
 wire \MuI._2427_ ;
 wire \MuI._2428_ ;
 wire \MuI._2429_ ;
 wire \MuI._2430_ ;
 wire \MuI._2431_ ;
 wire \MuI._2432_ ;
 wire \MuI._2433_ ;
 wire \MuI._2434_ ;
 wire \MuI._2435_ ;
 wire \MuI._2436_ ;
 wire \MuI._2437_ ;
 wire \MuI._2438_ ;
 wire \MuI._2439_ ;
 wire \MuI._2440_ ;
 wire \MuI._2441_ ;
 wire \MuI._2442_ ;
 wire \MuI._2443_ ;
 wire \MuI._2444_ ;
 wire \MuI._2445_ ;
 wire \MuI._2446_ ;
 wire \MuI._2447_ ;
 wire \MuI._2448_ ;
 wire \MuI._2449_ ;
 wire \MuI._2450_ ;
 wire \MuI._2451_ ;
 wire \MuI._2452_ ;
 wire \MuI._2453_ ;
 wire \MuI._2454_ ;
 wire \MuI._2455_ ;
 wire \MuI._2456_ ;
 wire \MuI._2457_ ;
 wire \MuI._2458_ ;
 wire \MuI._2459_ ;
 wire \MuI._2460_ ;
 wire \MuI._2461_ ;
 wire \MuI._2462_ ;
 wire \MuI._2463_ ;
 wire \MuI._2464_ ;
 wire \MuI._2465_ ;
 wire \MuI._2466_ ;
 wire \MuI._2467_ ;
 wire \MuI._2468_ ;
 wire \MuI._2469_ ;
 wire \MuI._2470_ ;
 wire \MuI._2471_ ;
 wire \MuI._2472_ ;
 wire \MuI._2473_ ;
 wire \MuI._2474_ ;
 wire \MuI._2475_ ;
 wire \MuI._2476_ ;
 wire \MuI._2477_ ;
 wire \MuI._2478_ ;
 wire \MuI._2479_ ;
 wire \MuI._2480_ ;
 wire \MuI._2481_ ;
 wire \MuI._2482_ ;
 wire \MuI._2483_ ;
 wire \MuI._2484_ ;
 wire \MuI._2485_ ;
 wire \MuI._2486_ ;
 wire \MuI._2487_ ;
 wire \MuI._2488_ ;
 wire \MuI._2489_ ;
 wire \MuI._2490_ ;
 wire \MuI._2491_ ;
 wire \MuI._2492_ ;
 wire \MuI._2493_ ;
 wire \MuI._2494_ ;
 wire \MuI._2495_ ;
 wire \MuI._2496_ ;
 wire \MuI._2497_ ;
 wire \MuI._2498_ ;
 wire \MuI._2499_ ;
 wire \MuI._2500_ ;
 wire \MuI._2501_ ;
 wire \MuI._2502_ ;
 wire \MuI._2503_ ;
 wire \MuI._2504_ ;
 wire \MuI._2505_ ;
 wire \MuI._2506_ ;
 wire \MuI._2507_ ;
 wire \MuI._2508_ ;
 wire \MuI._2509_ ;
 wire \MuI._2510_ ;
 wire \MuI._2511_ ;
 wire \MuI._2512_ ;
 wire \MuI._2513_ ;
 wire \MuI._2514_ ;
 wire \MuI._2515_ ;
 wire \MuI._2516_ ;
 wire \MuI._2517_ ;
 wire \MuI._2518_ ;
 wire \MuI._2519_ ;
 wire \MuI._2520_ ;
 wire \MuI._2521_ ;
 wire \MuI._2522_ ;
 wire \MuI._2523_ ;
 wire \MuI._2524_ ;
 wire \MuI._2525_ ;
 wire \MuI._2526_ ;
 wire \MuI._2527_ ;
 wire \MuI._2528_ ;
 wire \MuI._2529_ ;
 wire \MuI._2530_ ;
 wire \MuI._2531_ ;
 wire \MuI._2532_ ;
 wire \MuI._2533_ ;
 wire \MuI._2534_ ;
 wire \MuI._2535_ ;
 wire \MuI._2536_ ;
 wire \MuI._2537_ ;
 wire \MuI._2538_ ;
 wire \MuI._2539_ ;
 wire \MuI._2540_ ;
 wire \MuI._2541_ ;
 wire \MuI._2542_ ;
 wire \MuI._2543_ ;
 wire \MuI._2544_ ;
 wire \MuI._2545_ ;
 wire \MuI._2546_ ;
 wire \MuI._2547_ ;
 wire \MuI._2548_ ;
 wire \MuI._2549_ ;
 wire \MuI._2550_ ;
 wire \MuI._2551_ ;
 wire \MuI._2552_ ;
 wire \MuI._2553_ ;
 wire \MuI._2554_ ;
 wire \MuI._2555_ ;
 wire \MuI._2556_ ;
 wire \MuI._2557_ ;
 wire \MuI._2558_ ;
 wire \MuI._2559_ ;
 wire \MuI._2560_ ;
 wire \MuI._2561_ ;
 wire \MuI._2562_ ;
 wire \MuI._2563_ ;
 wire \MuI._2564_ ;
 wire \MuI._2565_ ;
 wire \MuI._2566_ ;
 wire \MuI._2567_ ;
 wire \MuI._2568_ ;
 wire \MuI._2569_ ;
 wire \MuI._2570_ ;
 wire \MuI._2571_ ;
 wire \MuI._2572_ ;
 wire \MuI._2573_ ;
 wire \MuI._2574_ ;
 wire \MuI._2575_ ;
 wire \MuI._2576_ ;
 wire \MuI._2577_ ;
 wire \MuI._2578_ ;
 wire \MuI._2579_ ;
 wire \MuI._2580_ ;
 wire \MuI._2581_ ;
 wire \MuI._2582_ ;
 wire \MuI._2583_ ;
 wire \MuI._2584_ ;
 wire \MuI._2585_ ;
 wire \MuI._2586_ ;
 wire \MuI._2587_ ;
 wire \MuI._2588_ ;
 wire \MuI._2589_ ;
 wire \MuI._2590_ ;
 wire \MuI._2591_ ;
 wire \MuI._2592_ ;
 wire \MuI._2593_ ;
 wire \MuI._2594_ ;
 wire \MuI._2595_ ;
 wire \MuI._2596_ ;
 wire \MuI._2597_ ;
 wire \MuI._2598_ ;
 wire \MuI._2599_ ;
 wire \MuI._2600_ ;
 wire \MuI._2601_ ;
 wire \MuI._2602_ ;
 wire \MuI._2603_ ;
 wire \MuI._2604_ ;
 wire \MuI._2605_ ;
 wire \MuI._2606_ ;
 wire \MuI._2607_ ;
 wire \MuI._2608_ ;
 wire \MuI._2609_ ;
 wire \MuI._2610_ ;
 wire \MuI._2611_ ;
 wire \MuI._2612_ ;
 wire \MuI._2613_ ;
 wire \MuI._2614_ ;
 wire \MuI._2615_ ;
 wire \MuI._2616_ ;
 wire \MuI._2617_ ;
 wire \MuI._2618_ ;
 wire \MuI._2619_ ;
 wire \MuI._2620_ ;
 wire \MuI._2621_ ;
 wire \MuI._2622_ ;
 wire \MuI._2623_ ;
 wire \MuI._2624_ ;
 wire \MuI._2625_ ;
 wire \MuI._2626_ ;
 wire \MuI._2627_ ;
 wire \MuI._2628_ ;
 wire \MuI._2629_ ;
 wire \MuI._2630_ ;
 wire \MuI._2631_ ;
 wire \MuI._2632_ ;
 wire \MuI._2633_ ;
 wire \MuI._2634_ ;
 wire \MuI._2635_ ;
 wire \MuI._2636_ ;
 wire \MuI._2637_ ;
 wire \MuI._2638_ ;
 wire \MuI._2639_ ;
 wire \MuI._2640_ ;
 wire \MuI._2641_ ;
 wire \MuI._2642_ ;
 wire \MuI._2643_ ;
 wire \MuI._2644_ ;
 wire \MuI._2645_ ;
 wire \MuI._2646_ ;
 wire \MuI._2647_ ;
 wire \MuI._2648_ ;
 wire \MuI._2649_ ;
 wire \MuI._2650_ ;
 wire \MuI._2651_ ;
 wire \MuI._2652_ ;
 wire \MuI._2653_ ;
 wire \MuI._2654_ ;
 wire \MuI._2655_ ;
 wire \MuI._2656_ ;
 wire \MuI._2657_ ;
 wire \MuI._2658_ ;
 wire \MuI._2659_ ;
 wire \MuI._2660_ ;
 wire \MuI._2661_ ;
 wire \MuI._2662_ ;
 wire \MuI._2663_ ;
 wire \MuI._2664_ ;
 wire \MuI._2665_ ;
 wire \MuI._2666_ ;
 wire \MuI._2667_ ;
 wire \MuI._2668_ ;
 wire \MuI._2669_ ;
 wire \MuI._2670_ ;
 wire \MuI._2671_ ;
 wire \MuI._2672_ ;
 wire \MuI._2673_ ;
 wire \MuI._2674_ ;
 wire \MuI._2675_ ;
 wire \MuI._2676_ ;
 wire \MuI._2677_ ;
 wire \MuI._2678_ ;
 wire \MuI._2679_ ;
 wire \MuI._2680_ ;
 wire \MuI._2681_ ;
 wire \MuI._2682_ ;
 wire \MuI._2683_ ;
 wire \MuI._2684_ ;
 wire \MuI._2685_ ;
 wire \MuI._2686_ ;
 wire \MuI._2687_ ;
 wire \MuI._2688_ ;
 wire \MuI._2689_ ;
 wire \MuI._2690_ ;
 wire \MuI._2691_ ;
 wire \MuI._2692_ ;
 wire \MuI._2693_ ;
 wire \MuI._2694_ ;
 wire \MuI._2695_ ;
 wire \MuI._2696_ ;
 wire \MuI._2697_ ;
 wire \MuI._2698_ ;
 wire \MuI._2699_ ;
 wire \MuI._2700_ ;
 wire \MuI._2701_ ;
 wire \MuI._2702_ ;
 wire \MuI._2703_ ;
 wire \MuI._2704_ ;
 wire \MuI._2705_ ;
 wire \MuI._2706_ ;
 wire \MuI._2707_ ;
 wire \MuI._2708_ ;
 wire \MuI._2709_ ;
 wire \MuI._2710_ ;
 wire \MuI._2711_ ;
 wire \MuI._2712_ ;
 wire \MuI._2713_ ;
 wire \MuI._2714_ ;
 wire \MuI._2715_ ;
 wire \MuI._2716_ ;
 wire \MuI._2717_ ;
 wire \MuI._2718_ ;
 wire \MuI._2719_ ;
 wire \MuI._2720_ ;
 wire \MuI._2721_ ;
 wire \MuI._2722_ ;
 wire \MuI._2723_ ;
 wire \MuI._2724_ ;
 wire \MuI._2725_ ;
 wire \MuI._2726_ ;
 wire \MuI._2727_ ;
 wire \MuI._2728_ ;
 wire \MuI._2729_ ;
 wire \MuI._2730_ ;
 wire \MuI._2731_ ;
 wire \MuI._2732_ ;
 wire \MuI._2733_ ;
 wire \MuI._2734_ ;
 wire \MuI._2735_ ;
 wire \MuI._2736_ ;
 wire \MuI._2737_ ;
 wire \MuI._2738_ ;
 wire \MuI._2739_ ;
 wire \MuI._2740_ ;
 wire \MuI._2741_ ;
 wire \MuI._2742_ ;
 wire \MuI._2743_ ;
 wire \MuI._2744_ ;
 wire \MuI._2745_ ;
 wire \MuI._2746_ ;
 wire \MuI._2747_ ;
 wire \MuI._2748_ ;
 wire \MuI._2749_ ;
 wire \MuI._2750_ ;
 wire \MuI._2751_ ;
 wire \MuI._2752_ ;
 wire \MuI._2753_ ;
 wire \MuI._2754_ ;
 wire \MuI._2755_ ;
 wire \MuI._2756_ ;
 wire \MuI._2757_ ;
 wire \MuI._2758_ ;
 wire \MuI._2759_ ;
 wire \MuI._2760_ ;
 wire \MuI._2761_ ;
 wire \MuI._2762_ ;
 wire \MuI._2763_ ;
 wire \MuI._2764_ ;
 wire \MuI._2765_ ;
 wire \MuI._2766_ ;
 wire \MuI._2767_ ;
 wire \MuI._2768_ ;
 wire \MuI._2769_ ;
 wire \MuI._2770_ ;
 wire \MuI._2771_ ;
 wire \MuI._2772_ ;
 wire \MuI._2773_ ;
 wire \MuI._2774_ ;
 wire \MuI._2775_ ;
 wire \MuI._2776_ ;
 wire \MuI._2777_ ;
 wire \MuI._2778_ ;
 wire \MuI._2779_ ;
 wire \MuI._2780_ ;
 wire \MuI._2781_ ;
 wire \MuI._2782_ ;
 wire \MuI._2783_ ;
 wire \MuI._2784_ ;
 wire \MuI._2785_ ;
 wire \MuI._2786_ ;
 wire \MuI._2787_ ;
 wire \MuI._2788_ ;
 wire \MuI._2789_ ;
 wire \MuI._2790_ ;
 wire \MuI._2791_ ;
 wire \MuI._2792_ ;
 wire \MuI._2793_ ;
 wire \MuI._2794_ ;
 wire \MuI._2795_ ;
 wire \MuI._2796_ ;
 wire \MuI._2797_ ;
 wire \MuI._2798_ ;
 wire \MuI._2799_ ;
 wire \MuI._2800_ ;
 wire \MuI._2801_ ;
 wire \MuI._2802_ ;
 wire \MuI._2803_ ;
 wire \MuI._2804_ ;
 wire \MuI._2805_ ;
 wire \MuI._2806_ ;
 wire \MuI._2807_ ;
 wire \MuI._2808_ ;
 wire \MuI._2809_ ;
 wire \MuI._2810_ ;
 wire \MuI._2811_ ;
 wire \MuI._2812_ ;
 wire \MuI._2813_ ;
 wire \MuI._2814_ ;
 wire \MuI._2815_ ;
 wire \MuI._2816_ ;
 wire \MuI._2817_ ;
 wire \MuI._2818_ ;
 wire \MuI._2819_ ;
 wire \MuI._2820_ ;
 wire \MuI._2821_ ;
 wire \MuI._2822_ ;
 wire \MuI._2823_ ;
 wire \MuI._2824_ ;
 wire \MuI._2825_ ;
 wire \MuI._2826_ ;
 wire \MuI._2827_ ;
 wire \MuI._2828_ ;
 wire \MuI._2829_ ;
 wire \MuI._2830_ ;
 wire \MuI._2831_ ;
 wire \MuI._2832_ ;
 wire \MuI._2833_ ;
 wire \MuI._2834_ ;
 wire \MuI._2835_ ;
 wire \MuI._2836_ ;
 wire \MuI._2837_ ;
 wire \MuI._2838_ ;
 wire \MuI._2839_ ;
 wire \MuI._2840_ ;
 wire \MuI._2841_ ;
 wire \MuI._2842_ ;
 wire \MuI._2843_ ;
 wire \MuI._2844_ ;
 wire \MuI._2845_ ;
 wire \MuI._2846_ ;
 wire \MuI._2847_ ;
 wire \MuI._2848_ ;
 wire \MuI._2849_ ;
 wire \MuI._2850_ ;
 wire \MuI._2851_ ;
 wire \MuI._2852_ ;
 wire \MuI._2853_ ;
 wire \MuI._2854_ ;
 wire \MuI._2855_ ;
 wire \MuI._2856_ ;
 wire \MuI._2857_ ;
 wire \MuI._2858_ ;
 wire \MuI._2859_ ;
 wire \MuI._2860_ ;
 wire \MuI._2861_ ;
 wire \MuI._2862_ ;
 wire \MuI._2863_ ;
 wire \MuI._2864_ ;
 wire \MuI._2865_ ;
 wire \MuI._2866_ ;
 wire \MuI._2867_ ;
 wire \MuI._2868_ ;
 wire \MuI._2869_ ;
 wire \MuI._2870_ ;
 wire \MuI._2871_ ;
 wire \MuI._2872_ ;
 wire \MuI._2873_ ;
 wire \MuI._2874_ ;
 wire \MuI._2875_ ;
 wire \MuI._2876_ ;
 wire \MuI._2877_ ;
 wire \MuI._2878_ ;
 wire \MuI._2879_ ;
 wire \MuI._2880_ ;
 wire \MuI._2881_ ;
 wire \MuI._2882_ ;
 wire \MuI._2883_ ;
 wire \MuI._2884_ ;
 wire \MuI._2885_ ;
 wire \MuI._2886_ ;
 wire \MuI._2887_ ;
 wire \MuI._2888_ ;
 wire \MuI._2889_ ;
 wire \MuI._2890_ ;
 wire \MuI._2891_ ;
 wire \MuI._2892_ ;
 wire \MuI._2893_ ;
 wire \MuI._2894_ ;
 wire \MuI._2895_ ;
 wire \MuI._2896_ ;
 wire \MuI._2897_ ;
 wire \MuI._2898_ ;
 wire \MuI._2899_ ;
 wire \MuI._2900_ ;
 wire \MuI._2901_ ;
 wire \MuI._2902_ ;
 wire \MuI._2903_ ;
 wire \MuI._2904_ ;
 wire \MuI._2905_ ;
 wire \MuI._2906_ ;
 wire \MuI._2907_ ;
 wire \MuI._2908_ ;
 wire \MuI._2909_ ;
 wire \MuI._2910_ ;
 wire \MuI._2911_ ;
 wire \MuI._2912_ ;
 wire \MuI._2913_ ;
 wire \MuI._2914_ ;
 wire \MuI._2915_ ;
 wire \MuI._2916_ ;
 wire \MuI._2917_ ;
 wire \MuI._2918_ ;
 wire \MuI._2919_ ;
 wire \MuI._2920_ ;
 wire \MuI._2921_ ;
 wire \MuI._2922_ ;
 wire \MuI._2923_ ;
 wire \MuI._2924_ ;
 wire \MuI._2925_ ;
 wire \MuI._2926_ ;
 wire \MuI._2927_ ;
 wire \MuI._2928_ ;
 wire \MuI._2929_ ;
 wire \MuI._2930_ ;
 wire \MuI._2931_ ;
 wire \MuI._2932_ ;
 wire \MuI._2933_ ;
 wire \MuI._2934_ ;
 wire \MuI._2935_ ;
 wire \MuI._2936_ ;
 wire \MuI._2937_ ;
 wire \MuI._2938_ ;
 wire \MuI._2939_ ;
 wire \MuI._2940_ ;
 wire \MuI._2941_ ;
 wire \MuI._2942_ ;
 wire \MuI._2943_ ;
 wire \MuI._2944_ ;
 wire \MuI._2945_ ;
 wire \MuI._2946_ ;
 wire \MuI._2947_ ;
 wire \MuI._2948_ ;
 wire \MuI._2949_ ;
 wire \MuI._2950_ ;
 wire \MuI._2951_ ;
 wire \MuI._2952_ ;
 wire \MuI._2953_ ;
 wire \MuI._2954_ ;
 wire \MuI._2955_ ;
 wire \MuI._2956_ ;
 wire \MuI._2957_ ;
 wire \MuI._2958_ ;
 wire \MuI._2959_ ;
 wire \MuI._2960_ ;
 wire \MuI._2961_ ;
 wire \MuI._2962_ ;
 wire \MuI._2963_ ;
 wire \MuI._2964_ ;
 wire \MuI._2965_ ;
 wire \MuI._2966_ ;
 wire \MuI._2967_ ;
 wire \MuI._2968_ ;
 wire \MuI._2969_ ;
 wire \MuI._2970_ ;
 wire \MuI._2971_ ;
 wire \MuI._2972_ ;
 wire \MuI._2973_ ;
 wire \MuI._2974_ ;
 wire \MuI._2975_ ;
 wire \MuI._2976_ ;
 wire \MuI._2977_ ;
 wire \MuI._2978_ ;
 wire \MuI._2979_ ;
 wire \MuI._2980_ ;
 wire \MuI._2981_ ;
 wire \MuI._2982_ ;
 wire \MuI._2983_ ;
 wire \MuI._2984_ ;
 wire \MuI._2985_ ;
 wire \MuI._2986_ ;
 wire \MuI._2987_ ;
 wire \MuI._2988_ ;
 wire \MuI._2989_ ;
 wire \MuI._2990_ ;
 wire \MuI._2991_ ;
 wire \MuI._2992_ ;
 wire \MuI._2993_ ;
 wire \MuI._2994_ ;
 wire \MuI._2995_ ;
 wire \MuI._2996_ ;
 wire \MuI._2997_ ;
 wire \MuI._2998_ ;
 wire \MuI._2999_ ;
 wire \MuI._3000_ ;
 wire \MuI._3001_ ;
 wire \MuI._3002_ ;
 wire \MuI._3003_ ;
 wire \MuI._3004_ ;
 wire \MuI._3005_ ;
 wire \MuI._3006_ ;
 wire \MuI._3007_ ;
 wire \MuI._3008_ ;
 wire \MuI._3009_ ;
 wire \MuI._3010_ ;
 wire \MuI._3011_ ;
 wire \MuI._3012_ ;
 wire \MuI._3013_ ;
 wire \MuI._3014_ ;
 wire \MuI._3015_ ;
 wire \MuI._3016_ ;
 wire \MuI._3017_ ;
 wire \MuI._3018_ ;
 wire \MuI._3019_ ;
 wire \MuI._3020_ ;
 wire \MuI._3021_ ;
 wire \MuI._3022_ ;
 wire \MuI._3023_ ;
 wire \MuI._3024_ ;
 wire \MuI._3025_ ;
 wire \MuI._3026_ ;
 wire \MuI._3027_ ;
 wire \MuI._3028_ ;
 wire \MuI._3029_ ;
 wire \MuI._3030_ ;
 wire \MuI._3031_ ;
 wire \MuI._3032_ ;
 wire \MuI._3033_ ;
 wire \MuI._3034_ ;
 wire \MuI._3035_ ;
 wire \MuI._3036_ ;
 wire \MuI._3037_ ;
 wire \MuI._3038_ ;
 wire \MuI._3039_ ;
 wire \MuI._3040_ ;
 wire \MuI._3041_ ;
 wire \MuI._3042_ ;
 wire \MuI._3043_ ;
 wire \MuI._3044_ ;
 wire \MuI._3045_ ;
 wire \MuI._3046_ ;
 wire \MuI._3047_ ;
 wire \MuI._3048_ ;
 wire \MuI._3049_ ;
 wire \MuI._3050_ ;
 wire \MuI._3051_ ;
 wire \MuI._3052_ ;
 wire \MuI._3053_ ;
 wire \MuI._3054_ ;
 wire \MuI._3055_ ;
 wire \MuI._3056_ ;
 wire \MuI._3057_ ;
 wire \MuI._3058_ ;
 wire \MuI._3059_ ;
 wire \MuI._3060_ ;
 wire \MuI._3061_ ;
 wire \MuI._3062_ ;
 wire \MuI._3063_ ;
 wire \MuI._3064_ ;
 wire \MuI._3065_ ;
 wire \MuI._3066_ ;
 wire \MuI._3067_ ;
 wire \MuI._3068_ ;
 wire \MuI._3069_ ;
 wire \MuI._3070_ ;
 wire \MuI._3071_ ;
 wire \MuI._3072_ ;
 wire \MuI._3073_ ;
 wire \MuI._3074_ ;
 wire \MuI._3075_ ;
 wire \MuI._3076_ ;
 wire \MuI._3077_ ;
 wire \MuI._3078_ ;
 wire \MuI._3079_ ;
 wire \MuI._3080_ ;
 wire \MuI._3081_ ;
 wire \MuI._3082_ ;
 wire \MuI._3083_ ;
 wire \MuI._3084_ ;
 wire \MuI._3085_ ;
 wire \MuI._3086_ ;
 wire \MuI._3087_ ;
 wire \MuI._3088_ ;
 wire \MuI._3089_ ;
 wire \MuI._3090_ ;
 wire \MuI._3091_ ;
 wire \MuI._3092_ ;
 wire \MuI._3093_ ;
 wire \MuI._3094_ ;
 wire \MuI._3095_ ;
 wire \MuI._3096_ ;
 wire \MuI._3097_ ;
 wire \MuI._3098_ ;
 wire \MuI._3099_ ;
 wire \MuI._3100_ ;
 wire \MuI._3101_ ;
 wire \MuI._3102_ ;
 wire \MuI._3103_ ;
 wire \MuI._3104_ ;
 wire \MuI._3105_ ;
 wire \MuI._3106_ ;
 wire \MuI._3107_ ;
 wire \MuI._3108_ ;
 wire \MuI._3109_ ;
 wire \MuI._3110_ ;
 wire \MuI._3111_ ;
 wire \MuI._3112_ ;
 wire \MuI._3113_ ;
 wire \MuI._3114_ ;
 wire \MuI._3115_ ;
 wire \MuI._3116_ ;
 wire \MuI._3117_ ;
 wire \MuI._3118_ ;
 wire \MuI._3119_ ;
 wire \MuI._3120_ ;
 wire \MuI._3121_ ;
 wire \MuI._3122_ ;
 wire \MuI._3123_ ;
 wire \MuI._3124_ ;
 wire \MuI._3125_ ;
 wire \MuI._3126_ ;
 wire \MuI._3127_ ;
 wire \MuI._3128_ ;
 wire \MuI._3129_ ;
 wire \MuI._3130_ ;
 wire \MuI._3131_ ;
 wire \MuI._3132_ ;
 wire \MuI._3133_ ;
 wire \MuI._3134_ ;
 wire \MuI._3135_ ;
 wire \MuI._3136_ ;
 wire \MuI._3137_ ;
 wire \MuI._3138_ ;
 wire \MuI._3139_ ;
 wire \MuI._3140_ ;
 wire \MuI._3141_ ;
 wire \MuI._3142_ ;
 wire \MuI._3143_ ;
 wire \MuI._3144_ ;
 wire \MuI._3145_ ;
 wire \MuI._3146_ ;
 wire \MuI._3147_ ;
 wire \MuI._3148_ ;
 wire \MuI._3149_ ;
 wire \MuI._3150_ ;
 wire \MuI._3151_ ;
 wire \MuI._3152_ ;
 wire \MuI._3153_ ;
 wire \MuI._3154_ ;
 wire \MuI._3155_ ;
 wire \MuI._3156_ ;
 wire \MuI._3157_ ;
 wire \MuI._3158_ ;
 wire \MuI._3159_ ;
 wire \MuI._3160_ ;
 wire \MuI._3161_ ;
 wire \MuI._3162_ ;
 wire \MuI._3163_ ;
 wire \MuI._3164_ ;
 wire \MuI._3165_ ;
 wire \MuI._3166_ ;
 wire \MuI._3167_ ;
 wire \MuI._3168_ ;
 wire \MuI._3169_ ;
 wire \MuI._3170_ ;
 wire \MuI._3171_ ;
 wire \MuI._3172_ ;
 wire \MuI._3173_ ;
 wire \MuI._3174_ ;
 wire \MuI._3175_ ;
 wire \MuI._3176_ ;
 wire \MuI._3177_ ;
 wire \MuI._3178_ ;
 wire \MuI._3179_ ;
 wire \MuI._3180_ ;
 wire \MuI._3181_ ;
 wire \MuI._3182_ ;
 wire \MuI._3183_ ;
 wire \MuI._3184_ ;
 wire \MuI._3185_ ;
 wire \MuI._3186_ ;
 wire \MuI._3187_ ;
 wire \MuI._3188_ ;
 wire \MuI._3189_ ;
 wire \MuI._3190_ ;
 wire \MuI._3191_ ;
 wire \MuI._3192_ ;
 wire \MuI._3193_ ;
 wire \MuI._3194_ ;
 wire \MuI._3195_ ;
 wire \MuI._3196_ ;
 wire \MuI._3197_ ;
 wire \MuI._3198_ ;
 wire \MuI._3199_ ;
 wire \MuI._3200_ ;
 wire \MuI._3201_ ;
 wire \MuI._3202_ ;
 wire \MuI._3203_ ;
 wire \MuI._3204_ ;
 wire \MuI._3205_ ;
 wire \MuI._3206_ ;
 wire \MuI._3207_ ;
 wire \MuI._3208_ ;
 wire \MuI._3209_ ;
 wire \MuI._3210_ ;
 wire \MuI._3211_ ;
 wire \MuI._3212_ ;
 wire \MuI._3213_ ;
 wire \MuI._3214_ ;
 wire \MuI._3215_ ;
 wire \MuI._3216_ ;
 wire \MuI._3217_ ;
 wire \MuI._3218_ ;
 wire \MuI._3219_ ;
 wire \MuI._3220_ ;
 wire \MuI._3221_ ;
 wire \MuI._3222_ ;
 wire \MuI._3223_ ;
 wire \MuI._3224_ ;
 wire \MuI._3225_ ;
 wire \MuI._3226_ ;
 wire \MuI._3227_ ;
 wire \MuI._3228_ ;
 wire \MuI._3229_ ;
 wire \MuI._3230_ ;
 wire \MuI._3231_ ;
 wire \MuI._3232_ ;
 wire \MuI._3233_ ;
 wire \MuI._3234_ ;
 wire \MuI._3235_ ;
 wire \MuI._3236_ ;
 wire \MuI._3237_ ;
 wire \MuI._3238_ ;
 wire \MuI._3239_ ;
 wire \MuI._3240_ ;
 wire \MuI._3241_ ;
 wire \MuI._3242_ ;
 wire \MuI._3243_ ;
 wire \MuI._3244_ ;
 wire \MuI._3245_ ;
 wire \MuI._3246_ ;
 wire \MuI._3247_ ;
 wire \MuI._3248_ ;
 wire \MuI._3249_ ;
 wire \MuI._3250_ ;
 wire \MuI._3251_ ;
 wire \MuI._3252_ ;
 wire \MuI._3253_ ;
 wire \MuI._3254_ ;
 wire \MuI._3255_ ;
 wire \MuI._3256_ ;
 wire \MuI._3257_ ;
 wire \MuI._3258_ ;
 wire \MuI._3259_ ;
 wire \MuI._3260_ ;
 wire \MuI._3261_ ;
 wire \MuI._3262_ ;
 wire \MuI._3263_ ;
 wire \MuI._3264_ ;
 wire \MuI._3265_ ;
 wire \MuI._3266_ ;
 wire \MuI._3267_ ;
 wire \MuI._3268_ ;
 wire \MuI._3269_ ;
 wire \MuI._3270_ ;
 wire \MuI._3271_ ;
 wire \MuI._3272_ ;
 wire \MuI._3273_ ;
 wire \MuI._3274_ ;
 wire \MuI._3275_ ;
 wire \MuI._3276_ ;
 wire \MuI._3277_ ;
 wire \MuI._3278_ ;
 wire \MuI._3279_ ;
 wire \MuI._3280_ ;
 wire \MuI._3281_ ;
 wire \MuI._3282_ ;
 wire \MuI._3283_ ;
 wire \MuI._3284_ ;
 wire \MuI._3285_ ;
 wire \MuI._3286_ ;
 wire \MuI._3287_ ;
 wire \MuI._3288_ ;
 wire \MuI._3289_ ;
 wire \MuI._3290_ ;
 wire \MuI._3291_ ;
 wire \MuI._3292_ ;
 wire \MuI._3293_ ;
 wire \MuI._3294_ ;
 wire \MuI._3295_ ;
 wire \MuI._3296_ ;
 wire \MuI._3297_ ;
 wire \MuI._3298_ ;
 wire \MuI._3299_ ;
 wire \MuI._3300_ ;
 wire \MuI._3301_ ;
 wire \MuI._3302_ ;
 wire \MuI._3303_ ;
 wire \MuI._3304_ ;
 wire \MuI._3305_ ;
 wire \MuI._3306_ ;
 wire \MuI._3307_ ;
 wire \MuI._3308_ ;
 wire \MuI._3309_ ;
 wire \MuI._3310_ ;
 wire \MuI._3311_ ;
 wire \MuI._3312_ ;
 wire \MuI._3313_ ;
 wire \MuI._3314_ ;
 wire \MuI._3315_ ;
 wire \MuI._3316_ ;
 wire \MuI._3317_ ;
 wire \MuI._3318_ ;
 wire \MuI._3319_ ;
 wire \MuI._3320_ ;
 wire \MuI._3321_ ;
 wire \MuI._3322_ ;
 wire \MuI._3323_ ;
 wire \MuI._3324_ ;
 wire \MuI._3325_ ;
 wire \MuI._3326_ ;
 wire \MuI._3327_ ;
 wire \MuI._3328_ ;
 wire \MuI._3329_ ;
 wire \MuI._3330_ ;
 wire \MuI._3331_ ;
 wire \MuI._3332_ ;
 wire \MuI._3333_ ;
 wire \MuI._3334_ ;
 wire \MuI._3335_ ;
 wire \MuI._3336_ ;
 wire \MuI._3337_ ;
 wire \MuI._3338_ ;
 wire \MuI._3339_ ;
 wire \MuI._3340_ ;
 wire \MuI._3341_ ;
 wire \MuI._3342_ ;
 wire \MuI._3343_ ;
 wire \MuI._3344_ ;
 wire \MuI._3345_ ;
 wire \MuI._3346_ ;
 wire \MuI._3347_ ;
 wire \MuI._3348_ ;
 wire \MuI._3349_ ;
 wire \MuI._3350_ ;
 wire \MuI._3351_ ;
 wire \MuI._3352_ ;
 wire \MuI._3353_ ;
 wire \MuI._3354_ ;
 wire \MuI._3355_ ;
 wire \MuI._3356_ ;
 wire \MuI._3357_ ;
 wire \MuI._3358_ ;
 wire \MuI._3359_ ;
 wire \MuI._3360_ ;
 wire \MuI._3361_ ;
 wire \MuI._3362_ ;
 wire \MuI._3363_ ;
 wire \MuI._3364_ ;
 wire \MuI._3365_ ;
 wire \MuI._3366_ ;
 wire \MuI._3367_ ;
 wire \MuI._3368_ ;
 wire \MuI._3369_ ;
 wire \MuI._3370_ ;
 wire \MuI._3371_ ;
 wire \MuI._3372_ ;
 wire \MuI._3373_ ;
 wire \MuI._3374_ ;
 wire \MuI._3375_ ;
 wire \MuI._3376_ ;
 wire \MuI._3377_ ;
 wire \MuI._3378_ ;
 wire \MuI._3379_ ;
 wire \MuI._3380_ ;
 wire \MuI._3381_ ;
 wire \MuI._3382_ ;
 wire \MuI._3383_ ;
 wire \MuI._3384_ ;
 wire \MuI._3385_ ;
 wire \MuI._3386_ ;
 wire \MuI._3387_ ;
 wire \MuI._3388_ ;
 wire \MuI._3389_ ;
 wire \MuI._3390_ ;
 wire \MuI._3391_ ;
 wire \MuI._3392_ ;
 wire \MuI._3393_ ;
 wire \MuI._3394_ ;
 wire \MuI._3395_ ;
 wire \MuI._3396_ ;
 wire \MuI._3397_ ;
 wire \MuI._3398_ ;
 wire \MuI._3399_ ;
 wire \MuI._3400_ ;
 wire \MuI._3401_ ;
 wire \MuI._3402_ ;
 wire \MuI._3403_ ;
 wire \MuI._3404_ ;
 wire \MuI._3405_ ;
 wire \MuI._3406_ ;
 wire \MuI._3407_ ;
 wire \MuI._3408_ ;
 wire \MuI._3409_ ;
 wire \MuI._3410_ ;
 wire \MuI._3411_ ;
 wire \MuI._3412_ ;
 wire \MuI._3413_ ;
 wire \MuI._3414_ ;
 wire \MuI._3415_ ;
 wire \MuI._3416_ ;
 wire \MuI._3417_ ;
 wire \MuI._3418_ ;
 wire \MuI._3419_ ;
 wire \MuI._3420_ ;
 wire \MuI._3421_ ;
 wire \MuI._3422_ ;
 wire \MuI.a_operand[0] ;
 wire \MuI.a_operand[10] ;
 wire \MuI.a_operand[11] ;
 wire \MuI.a_operand[12] ;
 wire \MuI.a_operand[13] ;
 wire \MuI.a_operand[14] ;
 wire \MuI.a_operand[15] ;
 wire \MuI.a_operand[16] ;
 wire \MuI.a_operand[17] ;
 wire \MuI.a_operand[18] ;
 wire \MuI.a_operand[19] ;
 wire \MuI.a_operand[1] ;
 wire \MuI.a_operand[20] ;
 wire \MuI.a_operand[21] ;
 wire \MuI.a_operand[22] ;
 wire \MuI.a_operand[23] ;
 wire \MuI.a_operand[24] ;
 wire \MuI.a_operand[25] ;
 wire \MuI.a_operand[26] ;
 wire \MuI.a_operand[27] ;
 wire \MuI.a_operand[28] ;
 wire \MuI.a_operand[29] ;
 wire \MuI.a_operand[2] ;
 wire \MuI.a_operand[30] ;
 wire \MuI.a_operand[31] ;
 wire \MuI.a_operand[3] ;
 wire \MuI.a_operand[4] ;
 wire \MuI.a_operand[5] ;
 wire \MuI.a_operand[6] ;
 wire \MuI.a_operand[7] ;
 wire \MuI.a_operand[8] ;
 wire \MuI.a_operand[9] ;
 wire \MuI.b_operand[0] ;
 wire \MuI.b_operand[10] ;
 wire \MuI.b_operand[11] ;
 wire \MuI.b_operand[12] ;
 wire \MuI.b_operand[13] ;
 wire \MuI.b_operand[14] ;
 wire \MuI.b_operand[15] ;
 wire \MuI.b_operand[16] ;
 wire \MuI.b_operand[17] ;
 wire \MuI.b_operand[18] ;
 wire \MuI.b_operand[19] ;
 wire \MuI.b_operand[1] ;
 wire \MuI.b_operand[20] ;
 wire \MuI.b_operand[21] ;
 wire \MuI.b_operand[22] ;
 wire \MuI.b_operand[23] ;
 wire \MuI.b_operand[24] ;
 wire \MuI.b_operand[25] ;
 wire \MuI.b_operand[26] ;
 wire \MuI.b_operand[27] ;
 wire \MuI.b_operand[28] ;
 wire \MuI.b_operand[29] ;
 wire \MuI.b_operand[2] ;
 wire \MuI.b_operand[30] ;
 wire \MuI.b_operand[31] ;
 wire \MuI.b_operand[3] ;
 wire \MuI.b_operand[4] ;
 wire \MuI.b_operand[5] ;
 wire \MuI.b_operand[6] ;
 wire \MuI.b_operand[7] ;
 wire \MuI.b_operand[8] ;
 wire \MuI.b_operand[9] ;
 wire \MuI.result[0] ;
 wire \MuI.result[10] ;
 wire \MuI.result[11] ;
 wire \MuI.result[12] ;
 wire \MuI.result[13] ;
 wire \MuI.result[14] ;
 wire \MuI.result[15] ;
 wire \MuI.result[16] ;
 wire \MuI.result[17] ;
 wire \MuI.result[18] ;
 wire \MuI.result[19] ;
 wire \MuI.result[1] ;
 wire \MuI.result[20] ;
 wire \MuI.result[21] ;
 wire \MuI.result[22] ;
 wire \MuI.result[23] ;
 wire \MuI.result[24] ;
 wire \MuI.result[25] ;
 wire \MuI.result[26] ;
 wire \MuI.result[27] ;
 wire \MuI.result[28] ;
 wire \MuI.result[29] ;
 wire \MuI.result[2] ;
 wire \MuI.result[30] ;
 wire \MuI.result[31] ;
 wire \MuI.result[3] ;
 wire \MuI.result[4] ;
 wire \MuI.result[5] ;
 wire \MuI.result[6] ;
 wire \MuI.result[7] ;
 wire \MuI.result[8] ;
 wire \MuI.result[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;

 sky130_fd_sc_hd__inv_2 \AuI._0805_  (.A(net20),
    .Y(\AuI._0025_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0806_  (.A(net18),
    .Y(\AuI._0026_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0807_  (.A(net17),
    .Y(\AuI._0027_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._0808_  (.A1(net50),
    .A2(\AuI._0026_ ),
    .B1(net49),
    .B2(\AuI._0027_ ),
    .X(\AuI._0028_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0809_  (.A(\AuI._0025_ ),
    .B(net114),
    .Y(\AuI._0029_ ));
 sky130_fd_sc_hd__and2_1 \AuI._0810_  (.A(\AuI._0025_ ),
    .B(net114),
    .X(\AuI._0030_ ));
 sky130_fd_sc_hd__or2_2 \AuI._0811_  (.A(\AuI._0029_ ),
    .B(\AuI._0030_ ),
    .X(\AuI._0031_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._0812_  (.A(net51),
    .B(net19),
    .X(\AuI._0032_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._0813_  (.A1(net50),
    .A2(\AuI._0026_ ),
    .B1(\AuI._0031_ ),
    .C1(\AuI._0032_ ),
    .X(\AuI._0033_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._0814_  (.A(net51),
    .B(\AuI._0030_ ),
    .C_N(net19),
    .X(\AuI._0034_ ));
 sky130_fd_sc_hd__o221a_1 \AuI._0815_  (.A1(\AuI._0025_ ),
    .A2(net114),
    .B1(\AuI._0028_ ),
    .B2(\AuI._0033_ ),
    .C1(\AuI._0034_ ),
    .X(\AuI._0035_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0816_  (.A(net119),
    .Y(\AuI._0036_ ));
 sky130_fd_sc_hd__or2_1 \AuI._0817_  (.A(\AuI._0036_ ),
    .B(net13),
    .X(\AuI._0037_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0818_  (.A(net117),
    .Y(\AuI._0038_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0819_  (.A(net118),
    .Y(\AuI._0039_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._0820_  (.A1(\AuI._0038_ ),
    .A2(net15),
    .B1(\AuI._0039_ ),
    .B2(net14),
    .X(\AuI._0040_ ));
 sky130_fd_sc_hd__or2_1 \AuI._0821_  (.A(\AuI._0038_ ),
    .B(net15),
    .X(\AuI._0041_ ));
 sky130_fd_sc_hd__or2_1 \AuI._0822_  (.A(\AuI._0039_ ),
    .B(net14),
    .X(\AuI._0042_ ));
 sky130_fd_sc_hd__and3b_1 \AuI._0823_  (.A_N(\AuI._0040_ ),
    .B(\AuI._0041_ ),
    .C(\AuI._0042_ ),
    .X(\AuI._0043_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0824_  (.A(net44),
    .Y(\AuI._0044_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._0825_  (.A1(\AuI._0036_ ),
    .A2(net13),
    .B1(\AuI._0044_ ),
    .B2(net133),
    .X(\AuI._0045_ ));
 sky130_fd_sc_hd__a32o_1 \AuI._0826_  (.A1(\AuI._0037_ ),
    .A2(\AuI._0043_ ),
    .A3(\AuI._0045_ ),
    .B1(\AuI._0041_ ),
    .B2(\AuI._0040_ ),
    .X(\AuI._0046_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0827_  (.A_N(net123),
    .B(net107),
    .X(\AuI._0047_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0828_  (.A_N(net124),
    .B(net108),
    .X(\AuI._0048_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0829_  (.A(\AuI._0047_ ),
    .B(\AuI._0048_ ),
    .Y(\AuI._0049_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0830_  (.A(net108),
    .Y(\AuI._0050_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0831_  (.A(net109),
    .Y(\AuI._0051_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._0832_  (.A1(\AuI._0050_ ),
    .A2(net124),
    .B1(net125),
    .B2(\AuI._0051_ ),
    .X(\AuI._0052_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0833_  (.A(net66),
    .Y(\AuI._0053_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0834_  (.A(net107),
    .Y(\AuI._0054_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._0835_  (.A1(\AuI._0053_ ),
    .A2(net34),
    .B1(\AuI._0054_ ),
    .B2(net123),
    .X(\AuI._0055_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0836_  (.A1(\AuI._0049_ ),
    .A2(\AuI._0052_ ),
    .B1(\AuI._0055_ ),
    .Y(\AuI._0056_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0837_  (.A(net27),
    .Y(\AuI._0057_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0838_  (.A(net116),
    .B_N(net132),
    .X(\AuI._0058_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0839_  (.A_N(net115),
    .B(net37),
    .X(\AuI._0059_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0840_  (.A_N(net132),
    .B(net116),
    .X(\AuI._0060_ ));
 sky130_fd_sc_hd__a221o_1 \AuI._0841_  (.A1(net111),
    .A2(\AuI._0057_ ),
    .B1(\AuI._0058_ ),
    .B2(\AuI._0059_ ),
    .C1(\AuI._0060_ ),
    .X(\AuI._0061_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0842_  (.A(net126),
    .Y(\AuI._0062_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._0843_  (.A1(net110),
    .A2(\AuI._0062_ ),
    .B1(net111),
    .B2(\AuI._0057_ ),
    .X(\AuI._0063_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0844_  (.A_N(net125),
    .B(net109),
    .X(\AuI._0064_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI._0845_  (.A1(net110),
    .A2(\AuI._0062_ ),
    .B1(\AuI._0047_ ),
    .C1(\AuI._0048_ ),
    .D1(\AuI._0064_ ),
    .X(\AuI._0065_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI._0846_  (.A1(\AuI._0061_ ),
    .A2(\AuI._0063_ ),
    .B1(\AuI._0065_ ),
    .C1(\AuI._0052_ ),
    .D1(\AuI._0055_ ),
    .X(\AuI._0066_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0847_  (.A(net120),
    .Y(\AuI._0067_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0848_  (.A(net121),
    .Y(\AuI._0068_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._0849_  (.A1(\AuI._0067_ ),
    .A2(net11),
    .B1(\AuI._0068_ ),
    .B2(net10),
    .X(\AuI._0069_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0850_  (.A(net8),
    .Y(\AuI._0070_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0851_  (.A(net41),
    .Y(\AuI._0071_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0852_  (.A1_N(\AuI._0070_ ),
    .A2_N(net40),
    .B1(\AuI._0071_ ),
    .B2(net9),
    .X(\AuI._0072_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._0853_  (.A1(\AuI._0068_ ),
    .A2(net10),
    .B1(\AuI._0071_ ),
    .B2(net9),
    .X(\AuI._0073_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0854_  (.A(net7),
    .Y(\AuI._0074_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0855_  (.A_N(net11),
    .B(net120),
    .X(\AuI._0075_ ));
 sky130_fd_sc_hd__a221oi_1 \AuI._0856_  (.A1(\AuI._0070_ ),
    .A2(net40),
    .B1(net122),
    .B2(\AuI._0074_ ),
    .C1(\AuI._0075_ ),
    .Y(\AuI._0076_ ));
 sky130_fd_sc_hd__or4bb_1 \AuI._0857_  (.A(\AuI._0069_ ),
    .B(\AuI._0072_ ),
    .C_N(\AuI._0073_ ),
    .D_N(\AuI._0076_ ),
    .X(\AuI._0077_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0858_  (.A(net38),
    .Y(\AuI._0078_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0859_  (.A1_N(net122),
    .A2_N(\AuI._0074_ ),
    .B1(\AuI._0078_ ),
    .B2(net6),
    .X(\AuI._0079_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0860_  (.A(net35),
    .Y(\AuI._0080_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0861_  (.A1_N(\AuI._0053_ ),
    .A2_N(net34),
    .B1(\AuI._0080_ ),
    .B2(net106),
    .X(\AuI._0081_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0862_  (.A(net68),
    .Y(\AuI._0082_ ));
 sky130_fd_sc_hd__o22ai_1 \AuI._0863_  (.A1(\AuI._0078_ ),
    .A2(net6),
    .B1(\AuI._0082_ ),
    .B2(net36),
    .Y(\AuI._0083_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0864_  (.A1_N(\AuI._0080_ ),
    .A2_N(net106),
    .B1(\AuI._0082_ ),
    .B2(net36),
    .X(\AuI._0084_ ));
 sky130_fd_sc_hd__or4_1 \AuI._0865_  (.A(\AuI._0079_ ),
    .B(\AuI._0081_ ),
    .C(\AuI._0083_ ),
    .D(\AuI._0084_ ),
    .X(\AuI._0085_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._0866_  (.A1(\AuI._0056_ ),
    .A2(\AuI._0066_ ),
    .B1(\AuI._0077_ ),
    .C1(\AuI._0085_ ),
    .X(\AuI._0086_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._0867_  (.A1(\AuI._0078_ ),
    .A2(net6),
    .B1(\AuI._0082_ ),
    .B2(net36),
    .X(\AuI._0087_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0868_  (.A1(\AuI._0087_ ),
    .A2(\AuI._0084_ ),
    .B1(\AuI._0079_ ),
    .Y(\AuI._0088_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0869_  (.A1(\AuI._0072_ ),
    .A2(\AuI._0073_ ),
    .B1(\AuI._0069_ ),
    .Y(\AuI._0089_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._0870_  (.A1(\AuI._0077_ ),
    .A2(\AuI._0088_ ),
    .B1(\AuI._0089_ ),
    .B2(\AuI._0075_ ),
    .X(\AuI._0090_ ));
 sky130_fd_sc_hd__o21ba_1 \AuI._0871_  (.A1(\AuI._0044_ ),
    .A2(net133),
    .B1_N(\AuI._0045_ ),
    .X(\AuI._0091_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._0872_  (.A(\AuI._0037_ ),
    .B(\AuI._0043_ ),
    .C(\AuI._0091_ ),
    .Y(\AuI._0092_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0873_  (.A1(\AuI._0086_ ),
    .A2(\AuI._0090_ ),
    .B1(\AuI._0092_ ),
    .Y(\AuI._0093_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0874_  (.A1(net49),
    .A2(\AuI._0027_ ),
    .B1(\AuI._0033_ ),
    .Y(\AuI._0094_ ));
 sky130_fd_sc_hd__o211ai_1 \AuI._0875_  (.A1(\AuI._0046_ ),
    .A2(\AuI._0093_ ),
    .B1(\AuI._0028_ ),
    .C1(\AuI._0094_ ),
    .Y(\AuI._0095_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._0876_  (.A(net112),
    .B(net131),
    .X(\AuI._0096_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._0877_  (.A(net55),
    .B(net23),
    .X(\AuI._0097_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0878_  (.A(net54),
    .B_N(net22),
    .X(\AuI._0098_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0879_  (.A(net22),
    .B_N(net54),
    .X(\AuI._0099_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._0880_  (.A(\AuI._0098_ ),
    .B(\AuI._0099_ ),
    .Y(\AuI._0100_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._0881_  (.A(net21),
    .B(net113),
    .X(\AuI._0101_ ));
 sky130_fd_sc_hd__or4_1 \AuI._0882_  (.A(\AuI._0096_ ),
    .B(\AuI._0097_ ),
    .C(\AuI._0100_ ),
    .D(\AuI._0101_ ),
    .X(\AuI._0102_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0883_  (.A1(\AuI._0035_ ),
    .A2(\AuI._0095_ ),
    .B1(\AuI._0102_ ),
    .Y(\AuI._0103_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0884_  (.A(net21),
    .Y(\AuI._0104_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._0885_  (.A1(\AuI._0104_ ),
    .A2(net113),
    .B1(\AuI._0098_ ),
    .Y(\AuI._0105_ ));
 sky130_fd_sc_hd__and4bb_1 \AuI._0886_  (.A_N(\AuI._0096_ ),
    .B_N(\AuI._0097_ ),
    .C(\AuI._0099_ ),
    .D(\AuI._0105_ ),
    .X(\AuI._0106_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0887_  (.A(net56),
    .Y(\AuI._0107_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._0888_  (.A1(\AuI._0107_ ),
    .A2(net131),
    .B1(net23),
    .Y(\AuI._0108_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0889_  (.A1_N(\AuI._0108_ ),
    .A2_N(net55),
    .B1(net131),
    .B2(\AuI._0107_ ),
    .X(\AuI._0109_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._0890_  (.A(net57),
    .B(net129),
    .Y(\AuI._0110_ ));
 sky130_fd_sc_hd__o31a_1 \AuI._0891_  (.A1(\AuI._0103_ ),
    .A2(\AuI._0106_ ),
    .A3(\AuI._0109_ ),
    .B1(\AuI._0110_ ),
    .X(\AuI._0111_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0892_  (.A(net129),
    .Y(\AuI._0112_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0893_  (.A(net58),
    .B_N(net128),
    .X(\AuI._0113_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._0894_  (.A1(net57),
    .A2(\AuI._0112_ ),
    .B1(\AuI._0113_ ),
    .Y(\AuI._0114_ ));
 sky130_fd_sc_hd__and2_1 \AuI._0895_  (.A(net28),
    .B(net60),
    .X(\AuI._0115_ ));
 sky130_fd_sc_hd__nor2_2 \AuI._0896_  (.A(net28),
    .B(net60),
    .Y(\AuI._0116_ ));
 sky130_fd_sc_hd__or2_2 \AuI._0897_  (.A(\AuI._0115_ ),
    .B(\AuI._0116_ ),
    .X(\AuI._0117_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0898_  (.A(net128),
    .B_N(net58),
    .X(\AuI._0118_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._0899_  (.A1(\AuI._0111_ ),
    .A2(\AuI._0114_ ),
    .B1(\AuI._0117_ ),
    .C1(\AuI._0118_ ),
    .X(\AuI._0119_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0900_  (.A_N(net60),
    .B(net28),
    .X(\AuI._0120_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0901_  (.A(\AuI._0119_ ),
    .B(\AuI._0120_ ),
    .Y(\AuI._0121_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0902_  (.A(\AuI._0121_ ),
    .X(\AuI._0122_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0903_  (.A(\AuI._0122_ ),
    .X(\AuI._0123_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0904_  (.A(\AuI._0123_ ),
    .X(\AuI._0124_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0905_  (.A(\AuI._0124_ ),
    .X(\AuI._0125_ ));
 sky130_fd_sc_hd__buf_4 \AuI._0906_  (.A(\AuI._0125_ ),
    .X(\AuI._0126_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0907_  (.A0(net20),
    .A1(net114),
    .S(\AuI._0126_ ),
    .X(\AuI._0127_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0908_  (.A(\AuI._0127_ ),
    .X(\AuI.exp_a ));
 sky130_fd_sc_hd__o211ai_2 \AuI._0909_  (.A1(\AuI._0111_ ),
    .A2(\AuI._0114_ ),
    .B1(\AuI._0117_ ),
    .C1(\AuI._0118_ ),
    .Y(\AuI._0128_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0910_  (.A(net60),
    .B_N(net28),
    .X(\AuI._0129_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0911_  (.A(net113),
    .B(\AuI._0128_ ),
    .C(\AuI._0129_ ),
    .X(\AuI._0130_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._0912_  (.A1(\AuI._0128_ ),
    .A2(\AuI._0129_ ),
    .B1(\AuI._0104_ ),
    .Y(\AuI._0131_ ));
 sky130_fd_sc_hd__or2_1 \AuI._0913_  (.A(\AuI._0130_ ),
    .B(\AuI._0131_ ),
    .X(\AuI._0132_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0914_  (.A(\AuI._0132_ ),
    .X(\AuI.operand_a[24] ));
 sky130_fd_sc_hd__mux2_1 \AuI._0915_  (.A0(net22),
    .A1(net54),
    .S(\AuI._0121_ ),
    .X(\AuI._0133_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0916_  (.A(\AuI._0133_ ),
    .X(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__mux2_1 \AuI._0917_  (.A0(net23),
    .A1(net55),
    .S(\AuI._0126_ ),
    .X(\AuI._0134_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0918_  (.A(\AuI._0134_ ),
    .X(\AuI.operand_a[26] ));
 sky130_fd_sc_hd__mux2_1 \AuI._0919_  (.A0(net131),
    .A1(net56),
    .S(\AuI._0122_ ),
    .X(\AuI._0135_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0920_  (.A(\AuI._0135_ ),
    .X(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__mux2_1 \AuI._0921_  (.A0(net129),
    .A1(net57),
    .S(\AuI._0126_ ),
    .X(\AuI._0136_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0922_  (.A(\AuI._0136_ ),
    .X(\AuI.operand_a[28] ));
 sky130_fd_sc_hd__mux2_1 \AuI._0923_  (.A0(net26),
    .A1(net58),
    .S(\AuI._0122_ ),
    .X(\AuI._0137_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0924_  (.A(\AuI._0137_ ),
    .X(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__inv_2 \AuI._0925_  (.A(\AuI._0116_ ),
    .Y(\AuI.operand_a[30] ));
 sky130_fd_sc_hd__xor2_4 \AuI._0926_  (.A(\AuI.AddBar_Sub ),
    .B(net61),
    .X(\AuI._0138_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._0927_  (.A(net29),
    .B(\AuI._0138_ ),
    .Y(\AuI._0139_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0928_  (.A0(net5),
    .A1(net37),
    .S(\AuI._0125_ ),
    .X(\AuI._0140_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0929_  (.A1(\AuI._0128_ ),
    .A2(\AuI._0129_ ),
    .B1(net52),
    .X(\AuI._0141_ ));
 sky130_fd_sc_hd__or3_1 \AuI._0930_  (.A(net20),
    .B(\AuI._0119_ ),
    .C(\AuI._0120_ ),
    .X(\AuI._0142_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._0931_  (.A1(\AuI._0031_ ),
    .A2(\AuI._0141_ ),
    .A3(\AuI._0142_ ),
    .B1(\AuI._0101_ ),
    .X(\AuI._0143_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0932_  (.A1(\AuI._0128_ ),
    .A2(\AuI._0129_ ),
    .B1(net53),
    .X(\AuI._0144_ ));
 sky130_fd_sc_hd__or3_1 \AuI._0933_  (.A(net21),
    .B(\AuI._0119_ ),
    .C(\AuI._0120_ ),
    .X(\AuI._0145_ ));
 sky130_fd_sc_hd__a2bb2o_1 \AuI._0934_  (.A1_N(\AuI._0130_ ),
    .A2_N(\AuI._0131_ ),
    .B1(\AuI._0144_ ),
    .B2(\AuI._0145_ ),
    .X(\AuI._0146_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0935_  (.A1(\AuI._0143_ ),
    .A2(\AuI._0146_ ),
    .B1(\AuI._0100_ ),
    .X(\AuI._0147_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0936_  (.A0(net54),
    .A1(net22),
    .S(\AuI._0121_ ),
    .X(\AuI._0148_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0937_  (.A(\AuI._0148_ ),
    .B_N(\AuI.operand_a[25] ),
    .X(\AuI._0149_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0938_  (.A1(\AuI._0147_ ),
    .A2(\AuI._0149_ ),
    .B1(\AuI._0097_ ),
    .X(\AuI._0150_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._0939_  (.A(\AuI._0097_ ),
    .B(\AuI._0147_ ),
    .C(\AuI._0149_ ),
    .Y(\AuI._0151_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._0940_  (.A(\AuI._0150_ ),
    .B(\AuI._0151_ ),
    .Y(\AuI._0152_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0941_  (.A(\AuI._0152_ ),
    .X(\AuI._0153_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._0942_  (.A(\AuI._0113_ ),
    .B(\AuI._0118_ ),
    .Y(\AuI._0154_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0943_  (.A0(net55),
    .A1(net23),
    .S(\AuI._0121_ ),
    .X(\AuI._0155_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0944_  (.A(\AuI._0155_ ),
    .B_N(\AuI._0097_ ),
    .X(\AuI._0156_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0945_  (.A1(\AuI._0150_ ),
    .A2(\AuI._0156_ ),
    .B1(\AuI._0096_ ),
    .X(\AuI._0157_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0946_  (.A0(net56),
    .A1(net131),
    .S(\AuI._0122_ ),
    .X(\AuI._0158_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0947_  (.A(\AuI._0158_ ),
    .B_N(\AuI.operand_a[27] ),
    .X(\AuI._0159_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0948_  (.A0(net57),
    .A1(net25),
    .S(\AuI._0122_ ),
    .X(\AuI._0160_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._0949_  (.A_N(\AuI._0110_ ),
    .B(\AuI._0160_ ),
    .X(\AuI._0161_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._0950_  (.A1(\AuI._0110_ ),
    .A2(\AuI._0157_ ),
    .A3(\AuI._0159_ ),
    .B1(\AuI._0161_ ),
    .X(\AuI._0162_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._0951_  (.A(\AuI._0154_ ),
    .B(\AuI._0162_ ),
    .Y(\AuI._0163_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0952_  (.A(\AuI._0163_ ),
    .X(\AuI._0164_ ));
 sky130_fd_sc_hd__a311o_1 \AuI._0953_  (.A1(\AuI._0110_ ),
    .A2(\AuI._0157_ ),
    .A3(\AuI._0159_ ),
    .B1(\AuI._0161_ ),
    .C1(\AuI._0154_ ),
    .X(\AuI._0165_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0954_  (.A0(net58),
    .A1(net26),
    .S(\AuI._0122_ ),
    .X(\AuI._0166_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._0955_  (.A(\AuI._0166_ ),
    .B_N(\AuI.operand_a[29] ),
    .X(\AuI._0167_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._0956_  (.A1(\AuI._0165_ ),
    .A2(\AuI._0167_ ),
    .B1(\AuI._0117_ ),
    .X(\AuI._0168_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0957_  (.A(\AuI._0168_ ),
    .X(\AuI._0169_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0958_  (.A0(net119),
    .A1(net13),
    .S(\AuI._0123_ ),
    .X(\AuI._0170_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0959_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0170_ ),
    .X(\AuI._0171_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0960_  (.A0(net44),
    .A1(net12),
    .S(\AuI._0123_ ),
    .X(\AuI._0172_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0961_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0172_ ),
    .X(\AuI._0173_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0962_  (.A(\AuI._0029_ ),
    .B(\AuI._0030_ ),
    .Y(\AuI._0174_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0963_  (.A(\AuI._0174_ ),
    .X(\AuI._0175_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0964_  (.A(\AuI._0175_ ),
    .X(\AuI._0176_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0965_  (.A0(\AuI._0171_ ),
    .A1(\AuI._0173_ ),
    .S(\AuI._0176_ ),
    .X(\AuI._0177_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0966_  (.A(\AuI._0122_ ),
    .X(\AuI._0178_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0967_  (.A0(net47),
    .A1(net15),
    .S(\AuI._0178_ ),
    .X(\AuI._0179_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0968_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0179_ ),
    .X(\AuI._0180_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0969_  (.A0(net118),
    .A1(net14),
    .S(\AuI._0178_ ),
    .X(\AuI._0181_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0970_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0181_ ),
    .X(\AuI._0182_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0971_  (.A0(\AuI._0180_ ),
    .A1(\AuI._0182_ ),
    .S(\AuI._0176_ ),
    .X(\AuI._0183_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0972_  (.A0(net50),
    .A1(net18),
    .S(\AuI._0178_ ),
    .X(\AuI._0184_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0973_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0184_ ),
    .X(\AuI._0185_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0974_  (.A0(net49),
    .A1(net17),
    .S(\AuI._0178_ ),
    .X(\AuI._0186_ ));
 sky130_fd_sc_hd__and3_1 \AuI._0975_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0186_ ),
    .X(\AuI._0187_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0976_  (.A0(\AuI._0185_ ),
    .A1(\AuI._0187_ ),
    .S(\AuI._0175_ ),
    .X(\AuI._0188_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0977_  (.A(\AuI._0031_ ),
    .X(\AuI._0189_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._0978_  (.A(\AuI._0154_ ),
    .B(\AuI._0162_ ),
    .X(\AuI._0190_ ));
 sky130_fd_sc_hd__a21oi_2 \AuI._0979_  (.A1(\AuI._0165_ ),
    .A2(\AuI._0167_ ),
    .B1(\AuI._0117_ ),
    .Y(\AuI._0191_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0980_  (.A(\AuI._0190_ ),
    .B(\AuI._0191_ ),
    .Y(\AuI._0192_ ));
 sky130_fd_sc_hd__or4_1 \AuI._0981_  (.A(\AuI._0155_ ),
    .B(\AuI._0158_ ),
    .C(\AuI._0160_ ),
    .D(\AuI._0166_ ),
    .X(\AuI._0193_ ));
 sky130_fd_sc_hd__and2_1 \AuI._0982_  (.A(\AuI._0141_ ),
    .B(\AuI._0142_ ),
    .X(\AuI._0194_ ));
 sky130_fd_sc_hd__and2_1 \AuI._0983_  (.A(\AuI._0144_ ),
    .B(\AuI._0145_ ),
    .X(\AuI._0195_ ));
 sky130_fd_sc_hd__or4_1 \AuI._0984_  (.A(\AuI._0115_ ),
    .B(\AuI._0194_ ),
    .C(\AuI._0195_ ),
    .D(\AuI._0148_ ),
    .X(\AuI._0196_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._0985_  (.A(\AuI._0193_ ),
    .B(\AuI._0196_ ),
    .Y(\AuI._0197_ ));
 sky130_fd_sc_hd__inv_2 \AuI._0986_  (.A(\AuI._0197_ ),
    .Y(\AuI._0198_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0987_  (.A(\AuI._0163_ ),
    .X(\AuI._0199_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._0988_  (.A(\AuI._0168_ ),
    .X(\AuI._0200_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._0989_  (.A0(net51),
    .A1(net19),
    .S(\AuI._0123_ ),
    .X(\AuI._0201_ ));
 sky130_fd_sc_hd__and4_1 \AuI._0990_  (.A(\AuI._0175_ ),
    .B(\AuI._0199_ ),
    .C(\AuI._0200_ ),
    .D(\AuI._0201_ ),
    .X(\AuI._0202_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._0991_  (.A1(\AuI._0189_ ),
    .A2(\AuI._0192_ ),
    .A3(\AuI._0198_ ),
    .B1(\AuI._0202_ ),
    .X(\AuI._0203_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._0992_  (.A(\AuI._0031_ ),
    .B(\AuI._0101_ ),
    .C(\AuI._0194_ ),
    .Y(\AuI._0204_ ));
 sky130_fd_sc_hd__and2_2 \AuI._0993_  (.A(\AuI._0143_ ),
    .B(\AuI._0204_ ),
    .X(\AuI._0205_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._0994_  (.A(\AuI._0205_ ),
    .X(\AuI._0206_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._0995_  (.A(\AuI._0143_ ),
    .B(\AuI._0146_ ),
    .Y(\AuI._0207_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._0996_  (.A(\AuI._0100_ ),
    .B(\AuI._0207_ ),
    .Y(\AuI._0208_ ));
 sky130_fd_sc_hd__buf_2 \AuI._0997_  (.A(\AuI._0208_ ),
    .X(\AuI._0209_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._0998_  (.A0(\AuI._0177_ ),
    .A1(\AuI._0183_ ),
    .A2(\AuI._0188_ ),
    .A3(\AuI._0203_ ),
    .S0(\AuI._0206_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0210_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._0999_  (.A(\AuI._0096_ ),
    .B(\AuI._0150_ ),
    .C(\AuI._0156_ ),
    .Y(\AuI._0211_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1000_  (.A(\AuI._0157_ ),
    .B(\AuI._0211_ ),
    .Y(\AuI._0212_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1001_  (.A1(\AuI._0153_ ),
    .A2(\AuI._0210_ ),
    .B1(\AuI._0212_ ),
    .X(\AuI._0213_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1002_  (.A0(net41),
    .A1(net9),
    .S(\AuI._0178_ ),
    .X(\AuI._0214_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1003_  (.A(\AuI._0190_ ),
    .B(\AuI._0191_ ),
    .C_N(\AuI._0214_ ),
    .X(\AuI._0215_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1004_  (.A0(net40),
    .A1(net8),
    .S(\AuI._0178_ ),
    .X(\AuI._0216_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1005_  (.A(\AuI._0190_ ),
    .B(\AuI._0191_ ),
    .C_N(\AuI._0216_ ),
    .X(\AuI._0217_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1006_  (.A0(net120),
    .A1(net11),
    .S(\AuI._0178_ ),
    .X(\AuI._0218_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1007_  (.A(\AuI._0190_ ),
    .B(\AuI._0191_ ),
    .C_N(\AuI._0218_ ),
    .X(\AuI._0219_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1008_  (.A0(net121),
    .A1(net10),
    .S(\AuI._0178_ ),
    .X(\AuI._0220_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1009_  (.A(\AuI._0190_ ),
    .B(\AuI._0191_ ),
    .C_N(\AuI._0220_ ),
    .X(\AuI._0221_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1010_  (.A0(\AuI._0215_ ),
    .A1(\AuI._0217_ ),
    .A2(\AuI._0219_ ),
    .A3(\AuI._0221_ ),
    .S0(\AuI._0176_ ),
    .S1(\AuI._0206_ ),
    .X(\AuI._0222_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1011_  (.A(\AuI._0143_ ),
    .B(\AuI._0204_ ),
    .Y(\AuI._0223_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1012_  (.A0(net122),
    .A1(net7),
    .S(\AuI._0123_ ),
    .X(\AuI._0224_ ));
 sky130_fd_sc_hd__a31oi_1 \AuI._1013_  (.A1(\AuI._0199_ ),
    .A2(\AuI._0200_ ),
    .A3(\AuI._0224_ ),
    .B1(\AuI._0176_ ),
    .Y(\AuI._0225_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1014_  (.A0(net38),
    .A1(net6),
    .S(\AuI._0123_ ),
    .X(\AuI._0226_ ));
 sky130_fd_sc_hd__a31oi_1 \AuI._1015_  (.A1(\AuI._0199_ ),
    .A2(\AuI._0200_ ),
    .A3(\AuI._0226_ ),
    .B1(\AuI._0189_ ),
    .Y(\AuI._0227_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1016_  (.A0(net67),
    .A1(net35),
    .S(\AuI._0122_ ),
    .X(\AuI._0228_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1017_  (.A0(net68),
    .A1(net36),
    .S(\AuI._0122_ ),
    .X(\AuI._0229_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1018_  (.A0(\AuI._0228_ ),
    .A1(\AuI._0229_ ),
    .S(\AuI._0031_ ),
    .X(\AuI._0230_ ));
 sky130_fd_sc_hd__or4b_1 \AuI._1019_  (.A(\AuI._0205_ ),
    .B(\AuI._0190_ ),
    .C(\AuI._0191_ ),
    .D_N(\AuI._0230_ ),
    .X(\AuI._0231_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1020_  (.A(\AuI._0207_ ),
    .B_N(\AuI._0100_ ),
    .X(\AuI._0232_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1021_  (.A(\AuI._0147_ ),
    .B(\AuI._0232_ ),
    .Y(\AuI._0233_ ));
 sky130_fd_sc_hd__o311a_1 \AuI._1022_  (.A1(\AuI._0223_ ),
    .A2(\AuI._0225_ ),
    .A3(\AuI._0227_ ),
    .B1(\AuI._0231_ ),
    .C1(\AuI._0233_ ),
    .X(\AuI._0234_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1023_  (.A1(\AuI._0209_ ),
    .A2(\AuI._0222_ ),
    .B1(\AuI._0234_ ),
    .C1(\AuI._0152_ ),
    .X(\AuI._0235_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1024_  (.A(\AuI._0192_ ),
    .X(\AuI._0236_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1025_  (.A0(net107),
    .A1(net33),
    .S(\AuI._0178_ ),
    .X(\AuI._0237_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1026_  (.A0(net66),
    .A1(net34),
    .S(\AuI._0122_ ),
    .X(\AuI._0238_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1027_  (.A0(\AuI._0237_ ),
    .A1(\AuI._0238_ ),
    .S(\AuI._0031_ ),
    .X(\AuI._0239_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1028_  (.A0(net108),
    .A1(net124),
    .A2(net109),
    .A3(net125),
    .S0(\AuI._0123_ ),
    .S1(\AuI._0175_ ),
    .X(\AuI._0240_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1029_  (.A0(\AuI._0239_ ),
    .A1(\AuI._0240_ ),
    .S(\AuI._0223_ ),
    .X(\AuI._0241_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1030_  (.A0(net116),
    .A1(net16),
    .A2(net37),
    .A3(net5),
    .S0(\AuI._0123_ ),
    .S1(\AuI._0175_ ),
    .X(\AuI._0242_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1031_  (.A0(net110),
    .A1(net30),
    .A2(net59),
    .A3(net27),
    .S0(\AuI._0123_ ),
    .S1(\AuI._0174_ ),
    .X(\AuI._0243_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1032_  (.A0(\AuI._0242_ ),
    .A1(\AuI._0243_ ),
    .S(\AuI._0205_ ),
    .X(\AuI._0244_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1033_  (.A0(\AuI._0241_ ),
    .A1(\AuI._0244_ ),
    .S(\AuI._0233_ ),
    .X(\AuI._0245_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1034_  (.A(\AuI._0157_ ),
    .B(\AuI._0211_ ),
    .X(\AuI._0246_ ));
 sky130_fd_sc_hd__a31oi_1 \AuI._1035_  (.A1(\AuI._0153_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0245_ ),
    .B1(\AuI._0246_ ),
    .Y(\AuI._0247_ ));
 sky130_fd_sc_hd__and2_2 \AuI._1036_  (.A(\AuI._0157_ ),
    .B(\AuI._0159_ ),
    .X(\AuI._0248_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1037_  (.A(\AuI._0110_ ),
    .B(\AuI._0248_ ),
    .Y(\AuI._0249_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1038_  (.A1(\AuI._0235_ ),
    .A2(\AuI._0247_ ),
    .B1(\AuI._0249_ ),
    .Y(\AuI._0250_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1039_  (.A(\AuI._0213_ ),
    .B(\AuI._0250_ ),
    .X(\AuI._0251_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \AuI._1040_  (.A(\AuI._0251_ ),
    .X(\AuI._0252_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1041_  (.A(\AuI._0140_ ),
    .B(\AuI._0252_ ),
    .Y(\AuI._0253_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1042_  (.A(\AuI._0139_ ),
    .B(\AuI._0253_ ),
    .Y(\AuI._0254_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1043_  (.A(net29),
    .B(\AuI._0138_ ),
    .X(\AuI._0255_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1044_  (.A(\AuI._0255_ ),
    .X(\AuI._0256_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1045_  (.A(\AuI._0256_ ),
    .X(\AuI._0257_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1046_  (.A(\AuI._0257_ ),
    .X(\AuI._0258_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1047_  (.A(\AuI._0258_ ),
    .X(\AuI._0259_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1048_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0252_ ),
    .B1(\AuI._0140_ ),
    .Y(\AuI._0260_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1049_  (.A(\AuI._0254_ ),
    .B(\AuI._0260_ ),
    .Y(\AuI.pe.significand[0] ));
 sky130_fd_sc_hd__xor2_4 \AuI._1050_  (.A(\AuI._0110_ ),
    .B(\AuI._0248_ ),
    .X(\AuI._0261_ ));
 sky130_fd_sc_hd__and2_2 \AuI._1051_  (.A(\AuI._0150_ ),
    .B(\AuI._0151_ ),
    .X(\AuI._0262_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1052_  (.A(\AuI._0262_ ),
    .X(\AuI._0263_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1053_  (.A0(\AuI._0229_ ),
    .A1(\AuI._0226_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0264_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1054_  (.A(\AuI._0192_ ),
    .B(\AuI._0264_ ),
    .X(\AuI._0265_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1055_  (.A(\AuI._0199_ ),
    .B(\AuI._0200_ ),
    .C(\AuI._0224_ ),
    .X(\AuI._0266_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1056_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0216_ ),
    .X(\AuI._0267_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1057_  (.A0(\AuI._0266_ ),
    .A1(\AuI._0267_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0268_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1058_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0214_ ),
    .X(\AuI._0269_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1059_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0220_ ),
    .X(\AuI._0270_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1060_  (.A0(\AuI._0269_ ),
    .A1(\AuI._0270_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0271_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1061_  (.A(\AuI._0164_ ),
    .B(\AuI._0169_ ),
    .C(\AuI._0218_ ),
    .X(\AuI._0272_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1062_  (.A0(\AuI._0173_ ),
    .A1(\AuI._0272_ ),
    .S(\AuI._0176_ ),
    .X(\AuI._0273_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._1063_  (.A(\AuI._0206_ ),
    .X(\AuI._0274_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1064_  (.A0(\AuI._0265_ ),
    .A1(\AuI._0268_ ),
    .A2(\AuI._0271_ ),
    .A3(\AuI._0273_ ),
    .S0(\AuI._0274_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0275_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1065_  (.A(\AuI._0233_ ),
    .X(\AuI._0276_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1066_  (.A0(\AuI._0228_ ),
    .A1(\AuI._0238_ ),
    .S(\AuI._0175_ ),
    .X(\AuI._0277_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1067_  (.A0(net64),
    .A1(net124),
    .S(\AuI._0178_ ),
    .X(\AuI._0278_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1068_  (.A0(\AuI._0237_ ),
    .A1(\AuI._0278_ ),
    .S(\AuI._0175_ ),
    .X(\AuI._0279_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1069_  (.A(\AuI._0223_ ),
    .B(\AuI._0199_ ),
    .C(\AuI._0200_ ),
    .D(\AuI._0279_ ),
    .X(\AuI._0280_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1070_  (.A1(\AuI._0206_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0277_ ),
    .B1(\AuI._0280_ ),
    .X(\AuI._0281_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1071_  (.A0(net59),
    .A1(net27),
    .A2(net48),
    .A3(net16),
    .S0(\AuI._0123_ ),
    .S1(\AuI._0175_ ),
    .X(\AuI._0282_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1072_  (.A1(\AuI._0199_ ),
    .A2(\AuI._0200_ ),
    .A3(\AuI._0282_ ),
    .B1(\AuI._0205_ ),
    .X(\AuI._0283_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1073_  (.A0(net63),
    .A1(net62),
    .A2(net31),
    .A3(net30),
    .S0(\AuI._0174_ ),
    .S1(\AuI._0124_ ),
    .X(\AuI._0284_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1074_  (.A1(\AuI._0199_ ),
    .A2(\AuI._0200_ ),
    .A3(\AuI._0284_ ),
    .B1(\AuI._0223_ ),
    .X(\AuI._0285_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1075_  (.A1(\AuI._0283_ ),
    .A2(\AuI._0285_ ),
    .B1(\AuI._0208_ ),
    .X(\AuI._0286_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1076_  (.A1(\AuI._0276_ ),
    .A2(\AuI._0281_ ),
    .B1(\AuI._0286_ ),
    .C1(\AuI._0153_ ),
    .X(\AuI._0287_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._1077_  (.A(\AuI._0246_ ),
    .X(\AuI._0288_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1078_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0275_ ),
    .B1(\AuI._0287_ ),
    .C1(\AuI._0288_ ),
    .X(\AuI._0289_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1079_  (.A0(\AuI._0171_ ),
    .A1(\AuI._0182_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0290_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1080_  (.A0(\AuI._0180_ ),
    .A1(\AuI._0187_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0291_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1081_  (.A(\AuI._0199_ ),
    .B(\AuI._0200_ ),
    .C(\AuI._0201_ ),
    .X(\AuI._0292_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1082_  (.A0(\AuI._0185_ ),
    .A1(\AuI._0292_ ),
    .S(\AuI._0189_ ),
    .X(\AuI._0293_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1083_  (.A(\AuI._0176_ ),
    .B(\AuI._0192_ ),
    .C(\AuI._0198_ ),
    .X(\AuI._0294_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1084_  (.A0(\AuI._0290_ ),
    .A1(\AuI._0291_ ),
    .A2(\AuI._0293_ ),
    .A3(\AuI._0294_ ),
    .S0(\AuI._0274_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0295_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1085_  (.A1(\AuI._0153_ ),
    .A2(\AuI._0295_ ),
    .B1(\AuI._0212_ ),
    .X(\AuI._0296_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1086_  (.A(\AuI._0261_ ),
    .B(\AuI._0289_ ),
    .C(\AuI._0296_ ),
    .X(\AuI._0297_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1087_  (.A(\AuI._0252_ ),
    .B(\AuI._0297_ ),
    .Y(\AuI._0298_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1088_  (.A0(net16),
    .A1(net48),
    .S(\AuI._0124_ ),
    .X(\AuI._0299_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1089_  (.A(\AuI._0139_ ),
    .B(\AuI._0298_ ),
    .C_N(\AuI._0299_ ),
    .X(\AuI._0300_ ));
 sky130_fd_sc_hd__o21bai_1 \AuI._1090_  (.A1(\AuI._0139_ ),
    .A2(\AuI._0298_ ),
    .B1_N(\AuI._0299_ ),
    .Y(\AuI._0301_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1091_  (.A1(\AuI._0300_ ),
    .A2(\AuI._0301_ ),
    .B1(\AuI._0254_ ),
    .Y(\AuI._0302_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1092_  (.A(\AuI._0254_ ),
    .B(\AuI._0300_ ),
    .C(\AuI._0301_ ),
    .X(\AuI._0303_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1093_  (.A(\AuI._0302_ ),
    .B(\AuI._0303_ ),
    .Y(\AuI.pe.significand[1] ));
 sky130_fd_sc_hd__a32o_1 \AuI._1094_  (.A1(\AuI._0261_ ),
    .A2(\AuI._0289_ ),
    .A3(\AuI._0296_ ),
    .B1(\AuI._0213_ ),
    .B2(\AuI._0250_ ),
    .X(\AuI._0304_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1095_  (.A0(\AuI._0180_ ),
    .A1(\AuI._0182_ ),
    .A2(\AuI._0185_ ),
    .A3(\AuI._0187_ ),
    .S0(\AuI._0175_ ),
    .S1(\AuI._0205_ ),
    .X(\AuI._0305_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1096_  (.A(\AuI._0209_ ),
    .B(\AuI._0305_ ),
    .X(\AuI._0306_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1097_  (.A(\AuI._0223_ ),
    .X(\AuI._0307_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1098_  (.A1(\AuI._0307_ ),
    .A2(\AuI._0203_ ),
    .B1(\AuI._0276_ ),
    .X(\AuI._0308_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1099_  (.A1(\AuI._0153_ ),
    .A2(\AuI._0306_ ),
    .A3(\AuI._0308_ ),
    .B1(\AuI._0212_ ),
    .X(\AuI._0309_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1100_  (.A0(\AuI._0269_ ),
    .A1(\AuI._0267_ ),
    .S(\AuI._0176_ ),
    .X(\AuI._0310_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1101_  (.A0(\AuI._0272_ ),
    .A1(\AuI._0270_ ),
    .S(\AuI._0175_ ),
    .X(\AuI._0311_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1102_  (.A(\AuI._0225_ ),
    .B(\AuI._0227_ ),
    .Y(\AuI._0312_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1103_  (.A0(\AuI._0177_ ),
    .A1(\AuI._0310_ ),
    .A2(\AuI._0311_ ),
    .A3(\AuI._0312_ ),
    .S0(\AuI._0233_ ),
    .S1(\AuI._0307_ ),
    .X(\AuI._0313_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1104_  (.A0(\AuI._0240_ ),
    .A1(\AuI._0243_ ),
    .S(\AuI._0223_ ),
    .X(\AuI._0314_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1105_  (.A0(\AuI._0230_ ),
    .A1(\AuI._0239_ ),
    .S(\AuI._0223_ ),
    .X(\AuI._0315_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1106_  (.A0(\AuI._0314_ ),
    .A1(\AuI._0315_ ),
    .S(\AuI._0208_ ),
    .X(\AuI._0316_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1107_  (.A1(\AuI._0152_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0316_ ),
    .B1(\AuI._0246_ ),
    .X(\AuI._0317_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1108_  (.A1(\AuI._0262_ ),
    .A2(\AuI._0313_ ),
    .B1(\AuI._0317_ ),
    .X(\AuI._0318_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1109_  (.A(\AuI._0261_ ),
    .B(\AuI._0309_ ),
    .C(\AuI._0318_ ),
    .X(\AuI._0319_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1110_  (.A(\AuI._0319_ ),
    .X(\AuI._0320_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1111_  (.A(\AuI._0304_ ),
    .B(\AuI._0320_ ),
    .Y(\AuI._0321_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1112_  (.A1(\AuI._0304_ ),
    .A2(\AuI._0320_ ),
    .B1(\AuI._0321_ ),
    .C1(\AuI._0255_ ),
    .X(\AuI._0322_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1113_  (.A0(net27),
    .A1(net59),
    .S(\AuI._0124_ ),
    .X(\AuI._0323_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1114_  (.A(\AuI._0322_ ),
    .B(\AuI._0323_ ),
    .X(\AuI._0324_ ));
 sky130_fd_sc_hd__a21bo_1 \AuI._1115_  (.A1(\AuI._0254_ ),
    .A2(\AuI._0301_ ),
    .B1_N(\AuI._0300_ ),
    .X(\AuI._0325_ ));
 sky130_fd_sc_hd__and2_2 \AuI._1116_  (.A(\AuI._0324_ ),
    .B(\AuI._0325_ ),
    .X(\AuI._0326_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1117_  (.A(\AuI._0324_ ),
    .B(\AuI._0325_ ),
    .Y(\AuI._0327_ ));
 sky130_fd_sc_hd__nor2_4 \AuI._1118_  (.A(\AuI._0326_ ),
    .B(\AuI._0327_ ),
    .Y(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__and2_1 \AuI._1119_  (.A(\AuI._0322_ ),
    .B(\AuI._0323_ ),
    .X(\AuI._0328_ ));
 sky130_fd_sc_hd__nor2_2 \AuI._1120_  (.A(\AuI._0328_ ),
    .B(\AuI._0326_ ),
    .Y(\AuI._0329_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1121_  (.A(\AuI._0209_ ),
    .X(\AuI._0330_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1122_  (.A0(\AuI._0180_ ),
    .A1(\AuI._0185_ ),
    .A2(\AuI._0187_ ),
    .A3(\AuI._0292_ ),
    .S0(\AuI._0206_ ),
    .S1(\AuI._0189_ ),
    .X(\AuI._0331_ ));
 sky130_fd_sc_hd__a41o_1 \AuI._1123_  (.A1(\AuI._0176_ ),
    .A2(\AuI._0307_ ),
    .A3(\AuI._0236_ ),
    .A4(\AuI._0198_ ),
    .B1(\AuI._0233_ ),
    .X(\AuI._0332_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1124_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0331_ ),
    .B1(\AuI._0332_ ),
    .Y(\AuI._0333_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1125_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0333_ ),
    .B1(\AuI._0288_ ),
    .X(\AuI._0334_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1126_  (.A0(\AuI._0268_ ),
    .A1(\AuI._0271_ ),
    .A2(\AuI._0273_ ),
    .A3(\AuI._0290_ ),
    .S0(\AuI._0206_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0335_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1127_  (.A(\AuI._0206_ ),
    .B(\AuI._0192_ ),
    .C(\AuI._0264_ ),
    .X(\AuI._0336_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1128_  (.A(\AuI._0307_ ),
    .B(\AuI._0192_ ),
    .C(\AuI._0277_ ),
    .X(\AuI._0337_ ));
 sky130_fd_sc_hd__a41o_1 \AuI._1129_  (.A1(\AuI._0223_ ),
    .A2(\AuI._0199_ ),
    .A3(\AuI._0200_ ),
    .A4(\AuI._0284_ ),
    .B1(\AuI._0208_ ),
    .X(\AuI._0338_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1130_  (.A1(\AuI._0206_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0279_ ),
    .B1(\AuI._0338_ ),
    .X(\AuI._0339_ ));
 sky130_fd_sc_hd__o311a_1 \AuI._1131_  (.A1(\AuI._0233_ ),
    .A2(\AuI._0336_ ),
    .A3(\AuI._0337_ ),
    .B1(\AuI._0339_ ),
    .C1(\AuI._0153_ ),
    .X(\AuI._0340_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1132_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0335_ ),
    .B1(\AuI._0340_ ),
    .C1(\AuI._0246_ ),
    .X(\AuI._0341_ ));
 sky130_fd_sc_hd__or3b_2 \AuI._1133_  (.A(\AuI._0334_ ),
    .B(\AuI._0249_ ),
    .C_N(\AuI._0341_ ),
    .X(\AuI._0342_ ));
 sky130_fd_sc_hd__o21bai_1 \AuI._1134_  (.A1(\AuI._0304_ ),
    .A2(\AuI._0320_ ),
    .B1_N(\AuI._0342_ ),
    .Y(\AuI._0343_ ));
 sky130_fd_sc_hd__nor3b_2 \AuI._1135_  (.A(\AuI._0304_ ),
    .B(\AuI._0320_ ),
    .C_N(\AuI._0342_ ),
    .Y(\AuI._0344_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1136_  (.A(\AuI._0344_ ),
    .Y(\AuI._0345_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1137_  (.A0(net30),
    .A1(net62),
    .S(\AuI._0125_ ),
    .X(\AuI._0346_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1138_  (.A(\AuI._0256_ ),
    .B(\AuI._0343_ ),
    .C(\AuI._0345_ ),
    .D(\AuI._0346_ ),
    .X(\AuI._0347_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1139_  (.A1(\AuI._0256_ ),
    .A2(\AuI._0343_ ),
    .A3(\AuI._0345_ ),
    .B1(\AuI._0346_ ),
    .X(\AuI._0348_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1140_  (.A_N(\AuI._0347_ ),
    .B(\AuI._0348_ ),
    .X(\AuI._0349_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1141_  (.A(\AuI._0329_ ),
    .B(\AuI._0349_ ),
    .Y(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__mux4_1 \AuI._1142_  (.A0(\AuI._0177_ ),
    .A1(\AuI._0183_ ),
    .A2(\AuI._0310_ ),
    .A3(\AuI._0311_ ),
    .S0(\AuI._0274_ ),
    .S1(\AuI._0276_ ),
    .X(\AuI._0350_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1143_  (.A(\AuI._0263_ ),
    .B(\AuI._0350_ ),
    .Y(\AuI._0351_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1144_  (.A(\AuI._0274_ ),
    .B(\AuI._0312_ ),
    .Y(\AuI._0352_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1145_  (.A1(\AuI._0236_ ),
    .A2(\AuI._0241_ ),
    .B1(\AuI._0209_ ),
    .Y(\AuI._0353_ ));
 sky130_fd_sc_hd__a311o_1 \AuI._1146_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0352_ ),
    .A3(\AuI._0231_ ),
    .B1(\AuI._0353_ ),
    .C1(\AuI._0262_ ),
    .X(\AuI._0354_ ));
 sky130_fd_sc_hd__a311o_1 \AuI._1147_  (.A1(\AuI._0189_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0198_ ),
    .B1(\AuI._0202_ ),
    .C1(\AuI._0307_ ),
    .X(\AuI._0355_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1148_  (.A1(\AuI._0274_ ),
    .A2(\AuI._0188_ ),
    .B1(\AuI._0355_ ),
    .Y(\AuI._0356_ ));
 sky130_fd_sc_hd__o31a_1 \AuI._1149_  (.A1(\AuI._0262_ ),
    .A2(\AuI._0330_ ),
    .A3(\AuI._0356_ ),
    .B1(\AuI._0288_ ),
    .X(\AuI._0357_ ));
 sky130_fd_sc_hd__a311o_2 \AuI._1150_  (.A1(\AuI._0212_ ),
    .A2(\AuI._0351_ ),
    .A3(\AuI._0354_ ),
    .B1(\AuI._0357_ ),
    .C1(\AuI._0249_ ),
    .X(\AuI._0358_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1151_  (.A(\AuI._0344_ ),
    .B(\AuI._0358_ ),
    .X(\AuI._0359_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1152_  (.A(\AuI._0344_ ),
    .B(\AuI._0358_ ),
    .Y(\AuI._0360_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1153_  (.A0(net31),
    .A1(net63),
    .S(\AuI._0124_ ),
    .X(\AuI._0361_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1154_  (.A(\AuI._0256_ ),
    .B(\AuI._0359_ ),
    .C(\AuI._0360_ ),
    .D(\AuI._0361_ ),
    .X(\AuI._0362_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1155_  (.A1(\AuI._0256_ ),
    .A2(\AuI._0359_ ),
    .A3(\AuI._0360_ ),
    .B1(\AuI._0361_ ),
    .X(\AuI._0363_ ));
 sky130_fd_sc_hd__and2b_2 \AuI._1156_  (.A_N(\AuI._0362_ ),
    .B(\AuI._0363_ ),
    .X(\AuI._0364_ ));
 sky130_fd_sc_hd__o31a_2 \AuI._1157_  (.A1(\AuI._0328_ ),
    .A2(\AuI._0326_ ),
    .A3(\AuI._0347_ ),
    .B1(\AuI._0348_ ),
    .X(\AuI._0365_ ));
 sky130_fd_sc_hd__xor2_4 \AuI._1158_  (.A(\AuI._0364_ ),
    .B(\AuI._0365_ ),
    .X(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__a21o_1 \AuI._1159_  (.A1(\AuI._0364_ ),
    .A2(\AuI._0365_ ),
    .B1(\AuI._0362_ ),
    .X(\AuI._0366_ ));
 sky130_fd_sc_hd__and4bb_1 \AuI._1160_  (.A_N(\AuI._0304_ ),
    .B_N(\AuI._0320_ ),
    .C(\AuI._0342_ ),
    .D(\AuI._0358_ ),
    .X(\AuI._0367_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1161_  (.A(\AuI._0307_ ),
    .B(\AuI._0236_ ),
    .C(\AuI._0264_ ),
    .X(\AuI._0368_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1162_  (.A1(\AuI._0274_ ),
    .A2(\AuI._0268_ ),
    .B1(\AuI._0368_ ),
    .C1(\AuI._0276_ ),
    .X(\AuI._0369_ ));
 sky130_fd_sc_hd__o211ai_2 \AuI._1163_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0281_ ),
    .B1(\AuI._0369_ ),
    .C1(\AuI._0153_ ),
    .Y(\AuI._0370_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1164_  (.A0(\AuI._0271_ ),
    .A1(\AuI._0273_ ),
    .A2(\AuI._0290_ ),
    .A3(\AuI._0291_ ),
    .S0(\AuI._0206_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0371_ ));
 sky130_fd_sc_hd__a21oi_2 \AuI._1165_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0371_ ),
    .B1(\AuI._0288_ ),
    .Y(\AuI._0372_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1166_  (.A1(\AuI._0176_ ),
    .A2(\AuI._0236_ ),
    .A3(\AuI._0198_ ),
    .B1(\AuI._0307_ ),
    .X(\AuI._0373_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1167_  (.A1(\AuI._0274_ ),
    .A2(\AuI._0293_ ),
    .B1(\AuI._0373_ ),
    .Y(\AuI._0374_ ));
 sky130_fd_sc_hd__or3_4 \AuI._1168_  (.A(\AuI._0262_ ),
    .B(\AuI._0330_ ),
    .C(\AuI._0374_ ),
    .X(\AuI._0375_ ));
 sky130_fd_sc_hd__a221oi_4 \AuI._1169_  (.A1(\AuI._0370_ ),
    .A2(\AuI._0372_ ),
    .B1(\AuI._0375_ ),
    .B2(\AuI._0288_ ),
    .C1(\AuI._0249_ ),
    .Y(\AuI._0376_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1170_  (.A(\AuI._0367_ ),
    .B(\AuI._0376_ ),
    .Y(\AuI._0377_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1171_  (.A0(net32),
    .A1(net64),
    .S(\AuI._0124_ ),
    .X(\AuI._0378_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._1172_  (.A(\AuI._0256_ ),
    .B(\AuI._0377_ ),
    .C(\AuI._0378_ ),
    .Y(\AuI._0379_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1173_  (.A1(\AuI._0256_ ),
    .A2(\AuI._0377_ ),
    .B1(\AuI._0378_ ),
    .X(\AuI._0380_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1174_  (.A(\AuI._0379_ ),
    .B(\AuI._0380_ ),
    .Y(\AuI._0381_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1175_  (.A(\AuI._0366_ ),
    .B(\AuI._0381_ ),
    .Y(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__a221o_2 \AuI._1176_  (.A1(\AuI._0370_ ),
    .A2(\AuI._0372_ ),
    .B1(\AuI._0375_ ),
    .B2(\AuI._0288_ ),
    .C1(\AuI._0249_ ),
    .X(\AuI._0382_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1177_  (.A0(\AuI._0177_ ),
    .A1(\AuI._0188_ ),
    .A2(\AuI._0311_ ),
    .A3(\AuI._0183_ ),
    .S0(\AuI._0208_ ),
    .S1(\AuI._0307_ ),
    .X(\AuI._0383_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1178_  (.A(\AuI._0199_ ),
    .B(\AuI._0200_ ),
    .C(\AuI._0226_ ),
    .X(\AuI._0384_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1179_  (.A0(\AuI._0266_ ),
    .A1(\AuI._0384_ ),
    .A2(\AuI._0269_ ),
    .A3(\AuI._0267_ ),
    .S0(\AuI._0176_ ),
    .S1(\AuI._0206_ ),
    .X(\AuI._0385_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1180_  (.A1(\AuI._0236_ ),
    .A2(\AuI._0315_ ),
    .B1(\AuI._0208_ ),
    .X(\AuI._0386_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1181_  (.A1(\AuI._0276_ ),
    .A2(\AuI._0385_ ),
    .B1(\AuI._0386_ ),
    .C1(\AuI._0153_ ),
    .X(\AuI._0387_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1182_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0383_ ),
    .B1(\AuI._0387_ ),
    .C1(\AuI._0288_ ),
    .X(\AuI._0388_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1183_  (.A(\AuI._0153_ ),
    .X(\AuI._0389_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1184_  (.A(\AuI._0307_ ),
    .B(\AuI._0203_ ),
    .X(\AuI._0390_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1185_  (.A1(\AuI._0389_ ),
    .A2(\AuI._0276_ ),
    .A3(\AuI._0390_ ),
    .B1(\AuI._0212_ ),
    .X(\AuI._0391_ ));
 sky130_fd_sc_hd__nand3_4 \AuI._1186_  (.A(\AuI._0261_ ),
    .B(\AuI._0388_ ),
    .C(\AuI._0391_ ),
    .Y(\AuI._0392_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1187_  (.A1(\AuI._0367_ ),
    .A2(\AuI._0382_ ),
    .B1(\AuI._0392_ ),
    .X(\AuI._0393_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._1188_  (.A(\AuI._0367_ ),
    .B(\AuI._0382_ ),
    .C(\AuI._0392_ ),
    .Y(\AuI._0394_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1189_  (.A0(net33),
    .A1(net65),
    .S(\AuI._0124_ ),
    .X(\AuI._0395_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1190_  (.A(\AuI._0255_ ),
    .B(\AuI._0393_ ),
    .C(\AuI._0394_ ),
    .D(\AuI._0395_ ),
    .X(\AuI._0396_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1191_  (.A1(\AuI._0256_ ),
    .A2(\AuI._0393_ ),
    .A3(\AuI._0394_ ),
    .B1(\AuI._0395_ ),
    .X(\AuI._0397_ ));
 sky130_fd_sc_hd__nand2b_2 \AuI._1192_  (.A_N(\AuI._0396_ ),
    .B(\AuI._0397_ ),
    .Y(\AuI._0398_ ));
 sky130_fd_sc_hd__and4b_1 \AuI._1193_  (.A_N(\AuI._0362_ ),
    .B(\AuI._0363_ ),
    .C(\AuI._0379_ ),
    .D(\AuI._0380_ ),
    .X(\AuI._0399_ ));
 sky130_fd_sc_hd__o311ai_2 \AuI._1194_  (.A1(\AuI._0328_ ),
    .A2(\AuI._0326_ ),
    .A3(\AuI._0347_ ),
    .B1(\AuI._0348_ ),
    .C1(\AuI._0399_ ),
    .Y(\AuI._0400_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1195_  (.A(\AuI._0256_ ),
    .B(\AuI._0377_ ),
    .C(\AuI._0378_ ),
    .X(\AuI._0401_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1196_  (.A1(\AuI._0362_ ),
    .A2(\AuI._0401_ ),
    .B1(\AuI._0380_ ),
    .Y(\AuI._0402_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1197_  (.A(\AuI._0400_ ),
    .B(\AuI._0402_ ),
    .X(\AuI._0403_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1198_  (.A(\AuI._0398_ ),
    .B(\AuI._0403_ ),
    .X(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__o21bai_2 \AuI._1199_  (.A1(\AuI._0398_ ),
    .A2(\AuI._0403_ ),
    .B1_N(\AuI._0396_ ),
    .Y(\AuI._0404_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1200_  (.A0(\AuI._0268_ ),
    .A1(\AuI._0271_ ),
    .S(\AuI._0274_ ),
    .X(\AuI._0405_ ));
 sky130_fd_sc_hd__o31a_1 \AuI._1201_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0336_ ),
    .A3(\AuI._0337_ ),
    .B1(\AuI._0153_ ),
    .X(\AuI._0406_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1202_  (.A1(\AuI._0276_ ),
    .A2(\AuI._0405_ ),
    .B1(\AuI._0406_ ),
    .Y(\AuI._0407_ ));
 sky130_fd_sc_hd__mux4_1 \AuI._1203_  (.A0(\AuI._0273_ ),
    .A1(\AuI._0290_ ),
    .A2(\AuI._0291_ ),
    .A3(\AuI._0293_ ),
    .S0(\AuI._0274_ ),
    .S1(\AuI._0209_ ),
    .X(\AuI._0408_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1204_  (.A1(\AuI._0263_ ),
    .A2(\AuI._0408_ ),
    .B1(\AuI._0288_ ),
    .Y(\AuI._0409_ ));
 sky130_fd_sc_hd__or4b_1 \AuI._1205_  (.A(\AuI._0262_ ),
    .B(\AuI._0330_ ),
    .C(\AuI._0274_ ),
    .D_N(\AuI._0294_ ),
    .X(\AuI._0410_ ));
 sky130_fd_sc_hd__a221o_2 \AuI._1206_  (.A1(\AuI._0407_ ),
    .A2(\AuI._0409_ ),
    .B1(\AuI._0410_ ),
    .B2(\AuI._0288_ ),
    .C1(\AuI._0249_ ),
    .X(\AuI._0411_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1207_  (.A1(\AuI._0367_ ),
    .A2(\AuI._0382_ ),
    .A3(\AuI._0392_ ),
    .B1(\AuI._0411_ ),
    .X(\AuI._0412_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1208_  (.A(\AuI._0358_ ),
    .B(\AuI._0382_ ),
    .C(\AuI._0392_ ),
    .D(\AuI._0411_ ),
    .X(\AuI._0413_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1209_  (.A1(\AuI._0344_ ),
    .A2(\AuI._0413_ ),
    .B1(\AuI._0139_ ),
    .Y(\AuI._0414_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1210_  (.A0(net34),
    .A1(net66),
    .S(\AuI._0124_ ),
    .X(\AuI._0415_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1211_  (.A(\AuI._0412_ ),
    .B(\AuI._0414_ ),
    .C(\AuI._0415_ ),
    .X(\AuI._0416_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1212_  (.A1(\AuI._0412_ ),
    .A2(\AuI._0414_ ),
    .B1(\AuI._0415_ ),
    .Y(\AuI._0417_ ));
 sky130_fd_sc_hd__or2_2 \AuI._1213_  (.A(\AuI._0416_ ),
    .B(\AuI._0417_ ),
    .X(\AuI._0418_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1214_  (.A(\AuI._0404_ ),
    .B(\AuI._0418_ ),
    .Y(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__and2_1 \AuI._1215_  (.A(\AuI._0344_ ),
    .B(\AuI._0413_ ),
    .X(\AuI._0419_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1216_  (.A(\AuI._0419_ ),
    .X(\AuI._0420_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1217_  (.A(\AuI._0288_ ),
    .B(\AuI._0249_ ),
    .Y(\AuI._0421_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1218_  (.A(\AuI._0421_ ),
    .X(\AuI._0422_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1219_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0222_ ),
    .B1(\AuI._0234_ ),
    .Y(\AuI._0423_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1220_  (.A0(\AuI._0210_ ),
    .A1(\AuI._0423_ ),
    .S(\AuI._0389_ ),
    .X(\AuI._0424_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1221_  (.A(\AuI._0422_ ),
    .B(\AuI._0424_ ),
    .Y(\AuI._0425_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1222_  (.A(\AuI._0420_ ),
    .B(\AuI._0425_ ),
    .Y(\AuI._0426_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1223_  (.A1(\AuI._0420_ ),
    .A2(\AuI._0425_ ),
    .B1(\AuI._0426_ ),
    .C1(\AuI._0139_ ),
    .X(\AuI._0427_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1224_  (.A0(net35),
    .A1(net67),
    .S(\AuI._0124_ ),
    .X(\AuI._0428_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1225_  (.A(\AuI._0427_ ),
    .B(\AuI._0428_ ),
    .X(\AuI._0429_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1226_  (.A(\AuI._0396_ ),
    .B(\AuI._0416_ ),
    .Y(\AuI._0430_ ));
 sky130_fd_sc_hd__o32a_1 \AuI._1227_  (.A1(\AuI._0398_ ),
    .A2(\AuI._0402_ ),
    .A3(\AuI._0418_ ),
    .B1(\AuI._0430_ ),
    .B2(\AuI._0417_ ),
    .X(\AuI._0431_ ));
 sky130_fd_sc_hd__o31a_1 \AuI._1228_  (.A1(\AuI._0398_ ),
    .A2(\AuI._0400_ ),
    .A3(\AuI._0418_ ),
    .B1(\AuI._0431_ ),
    .X(\AuI._0432_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1229_  (.A(\AuI._0429_ ),
    .B(\AuI._0432_ ),
    .X(\AuI._0433_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1230_  (.A(\AuI._0429_ ),
    .B(\AuI._0432_ ),
    .Y(\AuI._0434_ ));
 sky130_fd_sc_hd__nor2_2 \AuI._1231_  (.A(\AuI._0433_ ),
    .B(\AuI._0434_ ),
    .Y(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__and2b_1 \AuI._1232_  (.A_N(\AuI._0427_ ),
    .B(\AuI._0428_ ),
    .X(\AuI._0435_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1233_  (.A(\AuI._0435_ ),
    .B(\AuI._0434_ ),
    .Y(\AuI._0436_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1234_  (.A(\AuI._0256_ ),
    .X(\AuI._0437_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1235_  (.A(\AuI._0263_ ),
    .X(\AuI._0438_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1236_  (.A0(\AuI._0275_ ),
    .A1(\AuI._0295_ ),
    .S(\AuI._0438_ ),
    .X(\AuI._0439_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1237_  (.A(\AuI._0422_ ),
    .B(\AuI._0439_ ),
    .Y(\AuI._0440_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1238_  (.A1(\AuI._0420_ ),
    .A2(\AuI._0425_ ),
    .B1(\AuI._0440_ ),
    .X(\AuI._0441_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1239_  (.A(\AuI._0425_ ),
    .B(\AuI._0440_ ),
    .X(\AuI._0442_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1240_  (.A(\AuI._0420_ ),
    .B(\AuI._0442_ ),
    .Y(\AuI._0443_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1241_  (.A0(net36),
    .A1(net68),
    .S(\AuI._0124_ ),
    .X(\AuI._0444_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1242_  (.A(\AuI._0437_ ),
    .B(\AuI._0441_ ),
    .C(\AuI._0443_ ),
    .D(\AuI._0444_ ),
    .X(\AuI._0445_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1243_  (.A1(\AuI._0437_ ),
    .A2(\AuI._0441_ ),
    .A3(\AuI._0443_ ),
    .B1(\AuI._0444_ ),
    .X(\AuI._0446_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1244_  (.A_N(\AuI._0445_ ),
    .B(\AuI._0446_ ),
    .X(\AuI._0447_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1245_  (.A(\AuI._0436_ ),
    .B(\AuI._0447_ ),
    .Y(\AuI.pe.significand[9] ));
 sky130_fd_sc_hd__and3_1 \AuI._1246_  (.A(\AuI._0344_ ),
    .B(\AuI._0413_ ),
    .C(\AuI._0442_ ),
    .X(\AuI._0448_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1247_  (.A(\AuI._0306_ ),
    .B(\AuI._0308_ ),
    .X(\AuI._0449_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1248_  (.A1(\AuI._0438_ ),
    .A2(\AuI._0313_ ),
    .B1(\AuI._0421_ ),
    .X(\AuI._0450_ ));
 sky130_fd_sc_hd__o21ai_4 \AuI._1249_  (.A1(\AuI._0389_ ),
    .A2(\AuI._0449_ ),
    .B1(\AuI._0450_ ),
    .Y(\AuI._0451_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1250_  (.A(\AuI._0448_ ),
    .B(\AuI._0451_ ),
    .X(\AuI._0452_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1251_  (.A(\AuI._0448_ ),
    .B(\AuI._0451_ ),
    .Y(\AuI._0453_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1252_  (.A0(net6),
    .A1(net38),
    .S(\AuI._0125_ ),
    .X(\AuI._0454_ ));
 sky130_fd_sc_hd__nand4_1 \AuI._1253_  (.A(\AuI._0437_ ),
    .B(\AuI._0452_ ),
    .C(\AuI._0453_ ),
    .D(\AuI._0454_ ),
    .Y(\AuI._0455_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1254_  (.A1(\AuI._0437_ ),
    .A2(\AuI._0452_ ),
    .A3(\AuI._0453_ ),
    .B1(\AuI._0454_ ),
    .X(\AuI._0456_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1255_  (.A(\AuI._0455_ ),
    .B(\AuI._0456_ ),
    .X(\AuI._0457_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1256_  (.A1(\AuI._0435_ ),
    .A2(\AuI._0445_ ),
    .B1(\AuI._0446_ ),
    .X(\AuI._0458_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1257_  (.A1(\AuI._0434_ ),
    .A2(\AuI._0447_ ),
    .B1(\AuI._0458_ ),
    .X(\AuI._0459_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1258_  (.A(\AuI._0457_ ),
    .B(\AuI._0459_ ),
    .X(\AuI.pe.significand[10] ));
 sky130_fd_sc_hd__a21bo_1 \AuI._1259_  (.A1(\AuI._0457_ ),
    .A2(\AuI._0459_ ),
    .B1_N(\AuI._0455_ ),
    .X(\AuI._0460_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1260_  (.A(\AuI._0438_ ),
    .B(\AuI._0333_ ),
    .Y(\AuI._0461_ ));
 sky130_fd_sc_hd__o211a_2 \AuI._1261_  (.A1(\AuI._0438_ ),
    .A2(\AuI._0335_ ),
    .B1(\AuI._0421_ ),
    .C1(\AuI._0461_ ),
    .X(\AuI._0462_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1262_  (.A(\AuI._0462_ ),
    .Y(\AuI._0463_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1263_  (.A1(\AuI._0448_ ),
    .A2(\AuI._0451_ ),
    .B1(\AuI._0463_ ),
    .X(\AuI._0464_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1264_  (.A(\AuI._0442_ ),
    .B(\AuI._0451_ ),
    .C(\AuI._0463_ ),
    .X(\AuI._0465_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1265_  (.A(\AuI._0420_ ),
    .B(\AuI._0465_ ),
    .Y(\AuI._0466_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1266_  (.A0(net7),
    .A1(net122),
    .S(\AuI._0125_ ),
    .X(\AuI._0467_ ));
 sky130_fd_sc_hd__nand4_1 \AuI._1267_  (.A(\AuI._0437_ ),
    .B(\AuI._0464_ ),
    .C(\AuI._0466_ ),
    .D(\AuI._0467_ ),
    .Y(\AuI._0468_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1268_  (.A1(\AuI._0437_ ),
    .A2(\AuI._0464_ ),
    .A3(\AuI._0466_ ),
    .B1(\AuI._0467_ ),
    .X(\AuI._0469_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1269_  (.A(\AuI._0468_ ),
    .B(\AuI._0469_ ),
    .Y(\AuI._0470_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1270_  (.A(\AuI._0460_ ),
    .B(\AuI._0470_ ),
    .Y(\AuI.pe.significand[11] ));
 sky130_fd_sc_hd__nor2_1 \AuI._1271_  (.A(\AuI._0330_ ),
    .B(\AuI._0356_ ),
    .Y(\AuI._0471_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1272_  (.A(\AuI._0438_ ),
    .B(\AuI._0350_ ),
    .X(\AuI._0472_ ));
 sky130_fd_sc_hd__o211a_2 \AuI._1273_  (.A1(\AuI._0389_ ),
    .A2(\AuI._0471_ ),
    .B1(\AuI._0421_ ),
    .C1(\AuI._0472_ ),
    .X(\AuI._0473_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1274_  (.A(\AuI._0473_ ),
    .Y(\AuI._0474_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1275_  (.A1(\AuI._0420_ ),
    .A2(\AuI._0465_ ),
    .A3(\AuI._0474_ ),
    .B1(\AuI._0139_ ),
    .X(\AuI._0475_ ));
 sky130_fd_sc_hd__a21oi_4 \AuI._1276_  (.A1(\AuI._0466_ ),
    .A2(\AuI._0473_ ),
    .B1(\AuI._0475_ ),
    .Y(\AuI._0476_ ));
 sky130_fd_sc_hd__mux2_4 \AuI._1277_  (.A0(net8),
    .A1(net40),
    .S(\AuI._0125_ ),
    .X(\AuI._0477_ ));
 sky130_fd_sc_hd__xor2_4 \AuI._1278_  (.A(\AuI._0476_ ),
    .B(\AuI._0477_ ),
    .X(\AuI._0478_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1279_  (.A(\AuI._0455_ ),
    .B(\AuI._0456_ ),
    .C(\AuI._0468_ ),
    .D(\AuI._0469_ ),
    .X(\AuI._0479_ ));
 sky130_fd_sc_hd__nand3b_1 \AuI._1280_  (.A_N(\AuI._0429_ ),
    .B(\AuI._0447_ ),
    .C(\AuI._0479_ ),
    .Y(\AuI._0480_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1281_  (.A(\AuI._0455_ ),
    .B(\AuI._0468_ ),
    .Y(\AuI._0481_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._1282_  (.A1(\AuI._0458_ ),
    .A2(\AuI._0479_ ),
    .B1(\AuI._0481_ ),
    .B2(\AuI._0469_ ),
    .X(\AuI._0482_ ));
 sky130_fd_sc_hd__o21ba_2 \AuI._1283_  (.A1(\AuI._0432_ ),
    .A2(\AuI._0480_ ),
    .B1_N(\AuI._0482_ ),
    .X(\AuI._0483_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1284_  (.A(\AuI._0478_ ),
    .B(\AuI._0483_ ),
    .Y(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__and2_1 \AuI._1285_  (.A(\AuI._0476_ ),
    .B(\AuI._0477_ ),
    .X(\AuI._0484_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1286_  (.A_N(\AuI._0483_ ),
    .B(\AuI._0478_ ),
    .X(\AuI._0485_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1287_  (.A(\AuI._0420_ ),
    .B(\AuI._0465_ ),
    .C(\AuI._0474_ ),
    .X(\AuI._0486_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1288_  (.A(\AuI._0212_ ),
    .B(\AuI._0261_ ),
    .Y(\AuI._0487_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1289_  (.A(\AuI._0263_ ),
    .B(\AuI._0371_ ),
    .Y(\AuI._0488_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1290_  (.A1(\AuI._0330_ ),
    .A2(\AuI._0374_ ),
    .B1(\AuI._0263_ ),
    .X(\AuI._0489_ ));
 sky130_fd_sc_hd__or3_2 \AuI._1291_  (.A(\AuI._0487_ ),
    .B(\AuI._0488_ ),
    .C(\AuI._0489_ ),
    .X(\AuI._0490_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1292_  (.A(\AuI._0486_ ),
    .B(\AuI._0490_ ),
    .X(\AuI._0491_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1293_  (.A(\AuI._0486_ ),
    .B(\AuI._0490_ ),
    .Y(\AuI._0492_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1294_  (.A0(net9),
    .A1(net41),
    .S(\AuI._0125_ ),
    .X(\AuI._0493_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1295_  (.A(\AuI._0437_ ),
    .B(\AuI._0491_ ),
    .C(\AuI._0492_ ),
    .D(\AuI._0493_ ),
    .X(\AuI._0494_ ));
 sky130_fd_sc_hd__a31oi_2 \AuI._1296_  (.A1(\AuI._0257_ ),
    .A2(\AuI._0491_ ),
    .A3(\AuI._0492_ ),
    .B1(\AuI._0493_ ),
    .Y(\AuI._0495_ ));
 sky130_fd_sc_hd__o22ai_1 \AuI._1297_  (.A1(\AuI._0484_ ),
    .A2(\AuI._0485_ ),
    .B1(\AuI._0494_ ),
    .B2(\AuI._0495_ ),
    .Y(\AuI._0496_ ));
 sky130_fd_sc_hd__or4_1 \AuI._1298_  (.A(\AuI._0484_ ),
    .B(\AuI._0485_ ),
    .C(\AuI._0494_ ),
    .D(\AuI._0495_ ),
    .X(\AuI._0497_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1299_  (.A(\AuI._0496_ ),
    .B(\AuI._0497_ ),
    .Y(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__buf_2 \AuI._1300_  (.A(\AuI._0487_ ),
    .X(\AuI._0498_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1301_  (.A(\AuI._0438_ ),
    .B(\AuI._0383_ ),
    .Y(\AuI._0499_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1302_  (.A1(\AuI._0276_ ),
    .A2(\AuI._0390_ ),
    .B1(\AuI._0389_ ),
    .Y(\AuI._0500_ ));
 sky130_fd_sc_hd__or3_2 \AuI._1303_  (.A(\AuI._0498_ ),
    .B(\AuI._0499_ ),
    .C(\AuI._0500_ ),
    .X(\AuI._0501_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1304_  (.A1(\AuI._0486_ ),
    .A2(\AuI._0490_ ),
    .B1(\AuI._0501_ ),
    .X(\AuI._0502_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1305_  (.A(\AuI._0490_ ),
    .Y(\AuI._0503_ ));
 sky130_fd_sc_hd__nor3_1 \AuI._1306_  (.A(\AuI._0498_ ),
    .B(\AuI._0499_ ),
    .C(\AuI._0500_ ),
    .Y(\AuI._0504_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1307_  (.A(\AuI._0503_ ),
    .B(\AuI._0504_ ),
    .C_N(\AuI._0486_ ),
    .X(\AuI._0505_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1308_  (.A0(net10),
    .A1(net42),
    .S(\AuI._0125_ ),
    .X(\AuI._0506_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1309_  (.A(\AuI._0437_ ),
    .B(\AuI._0502_ ),
    .C(\AuI._0505_ ),
    .D(\AuI._0506_ ),
    .X(\AuI._0507_ ));
 sky130_fd_sc_hd__a31oi_2 \AuI._1310_  (.A1(\AuI._0437_ ),
    .A2(\AuI._0502_ ),
    .A3(\AuI._0505_ ),
    .B1(\AuI._0506_ ),
    .Y(\AuI._0508_ ));
 sky130_fd_sc_hd__nor2_2 \AuI._1311_  (.A(\AuI._0507_ ),
    .B(\AuI._0508_ ),
    .Y(\AuI._0509_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1312_  (.A(\AuI._0494_ ),
    .B(\AuI._0495_ ),
    .C_N(\AuI._0478_ ),
    .X(\AuI._0510_ ));
 sky130_fd_sc_hd__o21bai_1 \AuI._1313_  (.A1(\AuI._0484_ ),
    .A2(\AuI._0494_ ),
    .B1_N(\AuI._0495_ ),
    .Y(\AuI._0511_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1314_  (.A1(\AuI._0483_ ),
    .A2(\AuI._0510_ ),
    .B1(\AuI._0511_ ),
    .X(\AuI._0512_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1315_  (.A(\AuI._0509_ ),
    .B(\AuI._0512_ ),
    .Y(\AuI.pe.significand[14] ));
 sky130_fd_sc_hd__o21ba_1 \AuI._1316_  (.A1(\AuI._0508_ ),
    .A2(\AuI._0512_ ),
    .B1_N(\AuI._0507_ ),
    .X(\AuI._0513_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1317_  (.A1(\AuI._0276_ ),
    .A2(\AuI._0307_ ),
    .A3(\AuI._0294_ ),
    .B1(\AuI._0389_ ),
    .X(\AuI._0514_ ));
 sky130_fd_sc_hd__o211a_2 \AuI._1318_  (.A1(\AuI._0438_ ),
    .A2(\AuI._0408_ ),
    .B1(\AuI._0421_ ),
    .C1(\AuI._0514_ ),
    .X(\AuI._0515_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1319_  (.A(\AuI._0515_ ),
    .Y(\AuI._0516_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1320_  (.A1(\AuI._0486_ ),
    .A2(\AuI._0490_ ),
    .A3(\AuI._0501_ ),
    .B1(\AuI._0516_ ),
    .X(\AuI._0517_ ));
 sky130_fd_sc_hd__or4b_2 \AuI._1321_  (.A(\AuI._0503_ ),
    .B(\AuI._0504_ ),
    .C(\AuI._0515_ ),
    .D_N(\AuI._0486_ ),
    .X(\AuI._0518_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1322_  (.A0(net11),
    .A1(net120),
    .S(\AuI._0125_ ),
    .X(\AuI._0519_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1323_  (.A(\AuI._0437_ ),
    .B(\AuI._0517_ ),
    .C(\AuI._0518_ ),
    .D(\AuI._0519_ ),
    .X(\AuI._0520_ ));
 sky130_fd_sc_hd__a31oi_2 \AuI._1324_  (.A1(\AuI._0257_ ),
    .A2(\AuI._0517_ ),
    .A3(\AuI._0518_ ),
    .B1(\AuI._0519_ ),
    .Y(\AuI._0521_ ));
 sky130_fd_sc_hd__nor2_2 \AuI._1325_  (.A(\AuI._0520_ ),
    .B(\AuI._0521_ ),
    .Y(\AuI._0522_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1326_  (.A(\AuI._0513_ ),
    .B(\AuI._0522_ ),
    .Y(\AuI.pe.significand[15] ));
 sky130_fd_sc_hd__or3b_1 \AuI._1327_  (.A(\AuI._0498_ ),
    .B(\AuI._0438_ ),
    .C_N(\AuI._0210_ ),
    .X(\AuI._0523_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1328_  (.A(\AuI._0523_ ),
    .Y(\AuI._0524_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1329_  (.A(\AuI._0518_ ),
    .B(\AuI._0524_ ),
    .Y(\AuI._0525_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1330_  (.A1(\AuI._0518_ ),
    .A2(\AuI._0524_ ),
    .B1(\AuI._0525_ ),
    .C1(\AuI._0257_ ),
    .X(\AuI._0526_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1331_  (.A0(net12),
    .A1(net44),
    .S(\AuI._0125_ ),
    .X(\AuI._0527_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1332_  (.A(\AuI._0526_ ),
    .B(\AuI._0527_ ),
    .X(\AuI._0528_ ));
 sky130_fd_sc_hd__or4_1 \AuI._1333_  (.A(\AuI._0507_ ),
    .B(\AuI._0508_ ),
    .C(\AuI._0520_ ),
    .D(\AuI._0521_ ),
    .X(\AuI._0529_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1334_  (.A(\AuI._0510_ ),
    .B(\AuI._0529_ ),
    .Y(\AuI._0530_ ));
 sky130_fd_sc_hd__nor4_1 \AuI._1335_  (.A(\AuI._0432_ ),
    .B(\AuI._0480_ ),
    .C(\AuI._0510_ ),
    .D(\AuI._0529_ ),
    .Y(\AuI._0531_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1336_  (.A(\AuI._0507_ ),
    .B(\AuI._0520_ ),
    .Y(\AuI._0532_ ));
 sky130_fd_sc_hd__o22ai_1 \AuI._1337_  (.A1(\AuI._0521_ ),
    .A2(\AuI._0532_ ),
    .B1(\AuI._0529_ ),
    .B2(\AuI._0511_ ),
    .Y(\AuI._0533_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1338_  (.A1(\AuI._0482_ ),
    .A2(\AuI._0530_ ),
    .B1(\AuI._0531_ ),
    .C1(\AuI._0533_ ),
    .X(\AuI._0534_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1339_  (.A(\AuI._0528_ ),
    .B(\AuI._0534_ ),
    .X(\AuI.pe.significand[16] ));
 sky130_fd_sc_hd__nand2_1 \AuI._1340_  (.A(\AuI._0526_ ),
    .B(\AuI._0527_ ),
    .Y(\AuI._0535_ ));
 sky130_fd_sc_hd__a21bo_1 \AuI._1341_  (.A1(\AuI._0528_ ),
    .A2(\AuI._0534_ ),
    .B1_N(\AuI._0535_ ),
    .X(\AuI._0536_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1342_  (.A(\AuI._0389_ ),
    .B(\AuI._0295_ ),
    .C(\AuI._0422_ ),
    .X(\AuI._0537_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1343_  (.A1(\AuI._0518_ ),
    .A2(\AuI._0524_ ),
    .B1(\AuI._0537_ ),
    .Y(\AuI._0538_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1344_  (.A(\AuI._0486_ ),
    .B(\AuI._0490_ ),
    .C(\AuI._0501_ ),
    .D(\AuI._0516_ ),
    .X(\AuI._0539_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1345_  (.A(\AuI._0524_ ),
    .B(\AuI._0537_ ),
    .Y(\AuI._0540_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1346_  (.A1(\AuI._0539_ ),
    .A2(\AuI._0540_ ),
    .B1(\AuI._0139_ ),
    .Y(\AuI._0541_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1347_  (.A0(net13),
    .A1(net119),
    .S(\AuI._0126_ ),
    .X(\AuI._0542_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1348_  (.A(\AuI._0538_ ),
    .B(\AuI._0541_ ),
    .C(\AuI._0542_ ),
    .X(\AuI._0543_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1349_  (.A1(\AuI._0538_ ),
    .A2(\AuI._0541_ ),
    .B1(\AuI._0542_ ),
    .X(\AuI._0544_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1350_  (.A_N(\AuI._0543_ ),
    .B(\AuI._0544_ ),
    .X(\AuI._0545_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1351_  (.A(\AuI._0536_ ),
    .B(\AuI._0545_ ),
    .X(\AuI.pe.significand[17] ));
 sky130_fd_sc_hd__or3b_2 \AuI._1352_  (.A(\AuI._0498_ ),
    .B(\AuI._0438_ ),
    .C_N(\AuI._0449_ ),
    .X(\AuI._0546_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1353_  (.A1(\AuI._0539_ ),
    .A2(\AuI._0540_ ),
    .B1(\AuI._0546_ ),
    .Y(\AuI._0547_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1354_  (.A1(\AuI._0539_ ),
    .A2(\AuI._0540_ ),
    .A3(\AuI._0546_ ),
    .B1(\AuI._0139_ ),
    .X(\AuI._0548_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1355_  (.A(\AuI._0547_ ),
    .B(\AuI._0548_ ),
    .Y(\AuI._0549_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1356_  (.A0(net14),
    .A1(net46),
    .S(\AuI._0126_ ),
    .X(\AuI._0550_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1357_  (.A(\AuI._0549_ ),
    .B(\AuI._0550_ ),
    .X(\AuI._0551_ ));
 sky130_fd_sc_hd__a31oi_1 \AuI._1358_  (.A1(\AuI._0526_ ),
    .A2(\AuI._0527_ ),
    .A3(\AuI._0544_ ),
    .B1(\AuI._0543_ ),
    .Y(\AuI._0552_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1359_  (.A(\AuI._0552_ ),
    .Y(\AuI._0553_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1360_  (.A1(\AuI._0528_ ),
    .A2(\AuI._0534_ ),
    .A3(\AuI._0545_ ),
    .B1(\AuI._0553_ ),
    .X(\AuI._0554_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1361_  (.A(\AuI._0551_ ),
    .B(\AuI._0554_ ),
    .X(\AuI.pe.significand[18] ));
 sky130_fd_sc_hd__nand2_1 \AuI._1362_  (.A(\AuI._0549_ ),
    .B(\AuI._0550_ ),
    .Y(\AuI._0555_ ));
 sky130_fd_sc_hd__a21bo_1 \AuI._1363_  (.A1(\AuI._0551_ ),
    .A2(\AuI._0554_ ),
    .B1_N(\AuI._0555_ ),
    .X(\AuI._0556_ ));
 sky130_fd_sc_hd__or3_2 \AuI._1364_  (.A(\AuI._0438_ ),
    .B(\AuI._0333_ ),
    .C(\AuI._0498_ ),
    .X(\AuI._0557_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1365_  (.A1(\AuI._0539_ ),
    .A2(\AuI._0540_ ),
    .A3(\AuI._0546_ ),
    .B1(\AuI._0557_ ),
    .X(\AuI._0558_ ));
 sky130_fd_sc_hd__nand4_2 \AuI._1366_  (.A(\AuI._0539_ ),
    .B(\AuI._0540_ ),
    .C(\AuI._0546_ ),
    .D(\AuI._0557_ ),
    .Y(\AuI._0559_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1367_  (.A0(net15),
    .A1(net47),
    .S(\AuI._0126_ ),
    .X(\AuI._0560_ ));
 sky130_fd_sc_hd__nand4_1 \AuI._1368_  (.A(\AuI._0257_ ),
    .B(\AuI._0558_ ),
    .C(\AuI._0559_ ),
    .D(\AuI._0560_ ),
    .Y(\AuI._0561_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1369_  (.A1(\AuI._0257_ ),
    .A2(\AuI._0558_ ),
    .A3(\AuI._0559_ ),
    .B1(\AuI._0560_ ),
    .X(\AuI._0562_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1370_  (.A(\AuI._0561_ ),
    .B(\AuI._0562_ ),
    .X(\AuI._0563_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1371_  (.A(\AuI._0556_ ),
    .B(\AuI._0563_ ),
    .X(\AuI.pe.significand[19] ));
 sky130_fd_sc_hd__and3_1 \AuI._1372_  (.A(\AuI._0389_ ),
    .B(\AuI._0471_ ),
    .C(\AuI._0422_ ),
    .X(\AuI._0564_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1373_  (.A(\AuI._0559_ ),
    .B(\AuI._0564_ ),
    .X(\AuI._0565_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1374_  (.A0(net17),
    .A1(net49),
    .S(\AuI._0126_ ),
    .X(\AuI._0566_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1375_  (.A(\AuI._0257_ ),
    .B(\AuI._0565_ ),
    .C(\AuI._0566_ ),
    .X(\AuI._0567_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1376_  (.A1(\AuI._0257_ ),
    .A2(\AuI._0565_ ),
    .B1(\AuI._0566_ ),
    .Y(\AuI._0568_ ));
 sky130_fd_sc_hd__or2_2 \AuI._1377_  (.A(\AuI._0567_ ),
    .B(\AuI._0568_ ),
    .X(\AuI._0569_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1378_  (.A(\AuI._0528_ ),
    .B(\AuI._0545_ ),
    .C(\AuI._0551_ ),
    .D(\AuI._0563_ ),
    .X(\AuI._0570_ ));
 sky130_fd_sc_hd__and3b_1 \AuI._1379_  (.A_N(\AuI._0552_ ),
    .B(\AuI._0563_ ),
    .C(\AuI._0551_ ),
    .X(\AuI._0571_ ));
 sky130_fd_sc_hd__a21boi_1 \AuI._1380_  (.A1(\AuI._0555_ ),
    .A2(\AuI._0561_ ),
    .B1_N(\AuI._0562_ ),
    .Y(\AuI._0572_ ));
 sky130_fd_sc_hd__a211o_2 \AuI._1381_  (.A1(\AuI._0534_ ),
    .A2(\AuI._0570_ ),
    .B1(\AuI._0571_ ),
    .C1(\AuI._0572_ ),
    .X(\AuI._0573_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1382_  (.A(\AuI._0569_ ),
    .B(\AuI._0573_ ),
    .Y(\AuI.pe.significand[20] ));
 sky130_fd_sc_hd__nor2_1 \AuI._1383_  (.A(\AuI._0559_ ),
    .B(\AuI._0564_ ),
    .Y(\AuI._0574_ ));
 sky130_fd_sc_hd__or3_1 \AuI._1384_  (.A(\AuI._0375_ ),
    .B(\AuI._0498_ ),
    .C(\AuI._0574_ ),
    .X(\AuI._0575_ ));
 sky130_fd_sc_hd__o21ai_2 \AuI._1385_  (.A1(\AuI._0375_ ),
    .A2(\AuI._0498_ ),
    .B1(\AuI._0574_ ),
    .Y(\AuI._0576_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1386_  (.A0(net18),
    .A1(net50),
    .S(\AuI._0126_ ),
    .X(\AuI._0577_ ));
 sky130_fd_sc_hd__nand4_1 \AuI._1387_  (.A(\AuI._0257_ ),
    .B(\AuI._0575_ ),
    .C(\AuI._0576_ ),
    .D(\AuI._0577_ ),
    .Y(\AuI._0578_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1388_  (.A1(\AuI._0258_ ),
    .A2(\AuI._0575_ ),
    .A3(\AuI._0576_ ),
    .B1(\AuI._0577_ ),
    .X(\AuI._0579_ ));
 sky130_fd_sc_hd__nand2_2 \AuI._1389_  (.A(\AuI._0578_ ),
    .B(\AuI._0579_ ),
    .Y(\AuI._0580_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1390_  (.A(\AuI._0569_ ),
    .Y(\AuI._0581_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1391_  (.A1(\AuI._0581_ ),
    .A2(\AuI._0573_ ),
    .B1(\AuI._0567_ ),
    .X(\AuI._0582_ ));
 sky130_fd_sc_hd__xnor2_4 \AuI._1392_  (.A(\AuI._0580_ ),
    .B(\AuI._0582_ ),
    .Y(\AuI.pe.significand[21] ));
 sky130_fd_sc_hd__and4_1 \AuI._1393_  (.A(\AuI._0389_ ),
    .B(\AuI._0276_ ),
    .C(\AuI._0390_ ),
    .D(\AuI._0422_ ),
    .X(\AuI._0583_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1394_  (.A(\AuI._0576_ ),
    .B(\AuI._0583_ ),
    .Y(\AuI._0584_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1395_  (.A(\AuI._0576_ ),
    .B(\AuI._0583_ ),
    .X(\AuI._0585_ ));
 sky130_fd_sc_hd__mux2_2 \AuI._1396_  (.A0(net19),
    .A1(net51),
    .S(\AuI._0126_ ),
    .X(\AuI._0586_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1397_  (.A(\AuI._0258_ ),
    .B(\AuI._0584_ ),
    .C(\AuI._0585_ ),
    .D(\AuI._0586_ ),
    .X(\AuI._0587_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1398_  (.A1(\AuI._0258_ ),
    .A2(\AuI._0584_ ),
    .A3(\AuI._0585_ ),
    .B1(\AuI._0586_ ),
    .X(\AuI._0588_ ));
 sky130_fd_sc_hd__or2b_2 \AuI._1399_  (.A(\AuI._0587_ ),
    .B_N(\AuI._0588_ ),
    .X(\AuI._0589_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1400_  (.A(\AuI._0567_ ),
    .B_N(\AuI._0578_ ),
    .X(\AuI._0590_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1401_  (.A1(\AuI._0581_ ),
    .A2(\AuI._0573_ ),
    .B1(\AuI._0590_ ),
    .X(\AuI._0591_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1402_  (.A(\AuI._0579_ ),
    .B(\AuI._0591_ ),
    .Y(\AuI._0592_ ));
 sky130_fd_sc_hd__xor2_4 \AuI._1403_  (.A(\AuI._0589_ ),
    .B(\AuI._0592_ ),
    .X(\AuI.pe.significand[22] ));
 sky130_fd_sc_hd__a31o_1 \AuI._1404_  (.A1(\AuI._0579_ ),
    .A2(\AuI._0588_ ),
    .A3(\AuI._0591_ ),
    .B1(\AuI._0587_ ),
    .X(\AuI._0593_ ));
 sky130_fd_sc_hd__or4_1 \AuI._1405_  (.A(\AuI.operand_a[26] ),
    .B(\AuI.operand_a[27] ),
    .C(\AuI.operand_a[28] ),
    .D(\AuI.operand_a[29] ),
    .X(\AuI._0594_ ));
 sky130_fd_sc_hd__or4_1 \AuI._1406_  (.A(\AuI.operand_a[30] ),
    .B(\AuI.exp_a ),
    .C(\AuI.operand_a[24] ),
    .D(\AuI.operand_a[25] ),
    .X(\AuI._0595_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1407_  (.A(\AuI._0594_ ),
    .B(\AuI._0595_ ),
    .X(\AuI._0596_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1408_  (.A(\AuI._0576_ ),
    .B(\AuI._0583_ ),
    .Y(\AuI._0597_ ));
 sky130_fd_sc_hd__or2_2 \AuI._1409_  (.A(\AuI._0410_ ),
    .B(\AuI._0498_ ),
    .X(\AuI._0598_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI._1410_  (.A(\AuI._0139_ ),
    .X(\AuI._0599_ ));
 sky130_fd_sc_hd__a21oi_4 \AuI._1411_  (.A1(\AuI._0597_ ),
    .A2(\AuI._0598_ ),
    .B1(\AuI._0599_ ),
    .Y(\AuI.pe.significand[24] ));
 sky130_fd_sc_hd__o21a_1 \AuI._1412_  (.A1(\AuI._0597_ ),
    .A2(\AuI._0598_ ),
    .B1(\AuI.pe.significand[24] ),
    .X(\AuI._0600_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1413_  (.A(\AuI._0596_ ),
    .B(\AuI._0600_ ),
    .Y(\AuI._0601_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1414_  (.A(\AuI._0593_ ),
    .B(\AuI._0601_ ),
    .Y(\AuI.pe.significand[23] ));
 sky130_fd_sc_hd__nand3_1 \AuI._1415_  (.A(\AuI.exp_a ),
    .B(\AuI.operand_a[24] ),
    .C(\AuI.operand_a[25] ),
    .Y(\AuI._0602_ ));
 sky130_fd_sc_hd__inv_2 \AuI._1416_  (.A(\AuI._0602_ ),
    .Y(\AuI._0603_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1417_  (.A(\AuI.operand_a[26] ),
    .B(\AuI.operand_a[27] ),
    .C(\AuI._0603_ ),
    .X(\AuI._0604_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1418_  (.A(\AuI.operand_a[30] ),
    .B(\AuI.operand_a[28] ),
    .C(\AuI.operand_a[29] ),
    .D(\AuI._0604_ ),
    .X(\AuI._0605_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \AuI._1419_  (.A(\AuI._0605_ ),
    .X(\AuI.Exception ));
 sky130_fd_sc_hd__buf_2 \AuI._1420_  (.A(\AuI._0258_ ),
    .X(\AuI._0606_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1421_  (.A(\AuI._0140_ ),
    .B(\AuI._0252_ ),
    .X(\AuI._0607_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1422_  (.A(\AuI._0253_ ),
    .B(\AuI._0607_ ),
    .X(\AuI._0608_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1423_  (.A(\AuI._0261_ ),
    .B(\AuI._0289_ ),
    .C(\AuI._0296_ ),
    .D(\AuI._0299_ ),
    .X(\AuI._0609_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1424_  (.A1(\AuI._0261_ ),
    .A2(\AuI._0289_ ),
    .A3(\AuI._0296_ ),
    .B1(\AuI._0299_ ),
    .X(\AuI._0610_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1425_  (.A_N(\AuI._0609_ ),
    .B(\AuI._0610_ ),
    .X(\AuI._0611_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1426_  (.A(\AuI._0253_ ),
    .B(\AuI._0611_ ),
    .Y(\AuI._0612_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1427_  (.A_N(\AuI._0560_ ),
    .B(\AuI._0557_ ),
    .X(\AuI._0613_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1428_  (.A(\AuI._0546_ ),
    .B_N(\AuI._0550_ ),
    .X(\AuI._0614_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1429_  (.A(\AuI._0557_ ),
    .B_N(\AuI._0560_ ),
    .X(\AuI._0615_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1430_  (.A(\AuI._0560_ ),
    .B_N(\AuI._0557_ ),
    .X(\AuI._0616_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1431_  (.A(\AuI._0615_ ),
    .B(\AuI._0616_ ),
    .Y(\AuI._0617_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1432_  (.A1(\AuI._0389_ ),
    .A2(\AuI._0449_ ),
    .A3(\AuI._0422_ ),
    .B1(\AuI._0550_ ),
    .X(\AuI._0618_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1433_  (.A(\AuI._0614_ ),
    .B(\AuI._0618_ ),
    .Y(\AuI._0619_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1434_  (.A(\AuI._0617_ ),
    .B(\AuI._0619_ ),
    .X(\AuI._0620_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1435_  (.A(\AuI._0504_ ),
    .B(\AuI._0506_ ),
    .X(\AuI._0621_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1436_  (.A1(\AuI._0515_ ),
    .A2(\AuI._0519_ ),
    .B1(\AuI._0621_ ),
    .X(\AuI._0622_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1437_  (.A(\AuI._0503_ ),
    .B(\AuI._0493_ ),
    .X(\AuI._0623_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1438_  (.A(\AuI._0473_ ),
    .B(\AuI._0477_ ),
    .X(\AuI._0624_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1439_  (.A(\AuI._0515_ ),
    .B(\AuI._0519_ ),
    .X(\AuI._0625_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1440_  (.A(\AuI._0501_ ),
    .B(\AuI._0506_ ),
    .Y(\AuI._0626_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1441_  (.A(\AuI._0503_ ),
    .B(\AuI._0493_ ),
    .X(\AuI._0627_ ));
 sky130_fd_sc_hd__o2111a_1 \AuI._1442_  (.A1(\AuI._0623_ ),
    .A2(\AuI._0624_ ),
    .B1(\AuI._0625_ ),
    .C1(\AuI._0626_ ),
    .D1(\AuI._0627_ ),
    .X(\AuI._0628_ ));
 sky130_fd_sc_hd__a211oi_1 \AuI._1443_  (.A1(\AuI._0515_ ),
    .A2(\AuI._0519_ ),
    .B1(\AuI._0622_ ),
    .C1(\AuI._0628_ ),
    .Y(\AuI._0629_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1444_  (.A(\AuI._0503_ ),
    .B(\AuI._0493_ ),
    .Y(\AuI._0630_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1445_  (.A(\AuI._0625_ ),
    .B(\AuI._0626_ ),
    .Y(\AuI._0631_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1446_  (.A(\AuI._0473_ ),
    .B(\AuI._0477_ ),
    .Y(\AuI._0632_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1447_  (.A(\AuI._0624_ ),
    .B(\AuI._0632_ ),
    .Y(\AuI._0633_ ));
 sky130_fd_sc_hd__or4b_1 \AuI._1448_  (.A(\AuI._0630_ ),
    .B(\AuI._0631_ ),
    .C(\AuI._0623_ ),
    .D_N(\AuI._0633_ ),
    .X(\AuI._0634_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1449_  (.A(\AuI._0422_ ),
    .B(\AuI._0439_ ),
    .C(\AuI._0444_ ),
    .X(\AuI._0635_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1450_  (.A(\AuI._0422_ ),
    .B(\AuI._0424_ ),
    .C(\AuI._0428_ ),
    .X(\AuI._0636_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1451_  (.A1(\AuI._0422_ ),
    .A2(\AuI._0439_ ),
    .B1(\AuI._0444_ ),
    .X(\AuI._0637_ ));
 sky130_fd_sc_hd__xor2_2 \AuI._1452_  (.A(\AuI._0462_ ),
    .B(\AuI._0467_ ),
    .X(\AuI._0638_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1453_  (.A(\AuI._0451_ ),
    .B(\AuI._0454_ ),
    .Y(\AuI._0639_ ));
 sky130_fd_sc_hd__o2111a_1 \AuI._1454_  (.A1(\AuI._0635_ ),
    .A2(\AuI._0636_ ),
    .B1(\AuI._0637_ ),
    .C1(\AuI._0638_ ),
    .D1(\AuI._0639_ ),
    .X(\AuI._0640_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1455_  (.A_N(\AuI._0451_ ),
    .B(\AuI._0454_ ),
    .X(\AuI._0641_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1456_  (.A1(\AuI._0462_ ),
    .A2(\AuI._0467_ ),
    .B1(\AuI._0641_ ),
    .X(\AuI._0642_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1457_  (.A1(\AuI._0462_ ),
    .A2(\AuI._0467_ ),
    .B1(\AuI._0640_ ),
    .C1(\AuI._0642_ ),
    .X(\AuI._0643_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1458_  (.A(\AuI._0634_ ),
    .B_N(\AuI._0643_ ),
    .X(\AuI._0644_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1459_  (.A(\AuI._0411_ ),
    .B_N(\AuI._0415_ ),
    .X(\AuI._0645_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1460_  (.A(\AuI._0376_ ),
    .B(\AuI._0378_ ),
    .X(\AuI._0646_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1461_  (.A_N(\AuI._0358_ ),
    .B(\AuI._0361_ ),
    .X(\AuI._0647_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1462_  (.A(\AuI._0411_ ),
    .B(\AuI._0415_ ),
    .Y(\AuI._0648_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1463_  (.A(\AuI._0376_ ),
    .B(\AuI._0378_ ),
    .X(\AuI._0649_ ));
 sky130_fd_sc_hd__xnor2_2 \AuI._1464_  (.A(\AuI._0392_ ),
    .B(\AuI._0395_ ),
    .Y(\AuI._0650_ ));
 sky130_fd_sc_hd__o2111ai_4 \AuI._1465_  (.A1(\AuI._0646_ ),
    .A2(\AuI._0647_ ),
    .B1(\AuI._0648_ ),
    .C1(\AuI._0649_ ),
    .D1(\AuI._0650_ ),
    .Y(\AuI._0651_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1466_  (.A(\AuI._0346_ ),
    .B_N(\AuI._0342_ ),
    .X(\AuI._0652_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1467_  (.A(\AuI._0320_ ),
    .B(\AuI._0323_ ),
    .X(\AuI._0653_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1468_  (.A1(\AuI._0140_ ),
    .A2(\AuI._0252_ ),
    .A3(\AuI._0610_ ),
    .B1(\AuI._0609_ ),
    .X(\AuI._0654_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1469_  (.A_N(\AuI._0342_ ),
    .B(\AuI._0346_ ),
    .X(\AuI._0655_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1470_  (.A(\AuI._0320_ ),
    .B(\AuI._0323_ ),
    .X(\AuI._0656_ ));
 sky130_fd_sc_hd__a211o_1 \AuI._1471_  (.A1(\AuI._0653_ ),
    .A2(\AuI._0654_ ),
    .B1(\AuI._0655_ ),
    .C1(\AuI._0656_ ),
    .X(\AuI._0657_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1472_  (.A(\AuI._0358_ ),
    .B(\AuI._0361_ ),
    .Y(\AuI._0658_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1473_  (.A(\AuI._0382_ ),
    .B(\AuI._0378_ ),
    .Y(\AuI._0659_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1474_  (.A(\AuI._0650_ ),
    .B(\AuI._0658_ ),
    .C(\AuI._0659_ ),
    .D(\AuI._0648_ ),
    .X(\AuI._0660_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1475_  (.A_N(\AuI._0392_ ),
    .B(\AuI._0395_ ),
    .X(\AuI._0661_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1476_  (.A(\AuI._0415_ ),
    .B_N(\AuI._0411_ ),
    .X(\AuI._0662_ ));
 sky130_fd_sc_hd__a32oi_4 \AuI._1477_  (.A1(\AuI._0652_ ),
    .A2(\AuI._0657_ ),
    .A3(\AuI._0660_ ),
    .B1(\AuI._0661_ ),
    .B2(\AuI._0662_ ),
    .Y(\AuI._0663_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1478_  (.A(\AuI._0638_ ),
    .B(\AuI._0639_ ),
    .Y(\AuI._0664_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1479_  (.A1(\AuI._0422_ ),
    .A2(\AuI._0424_ ),
    .B1(\AuI._0428_ ),
    .Y(\AuI._0665_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1480_  (.A(\AuI._0636_ ),
    .B(\AuI._0665_ ),
    .X(\AuI._0666_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1481_  (.A_N(\AuI._0635_ ),
    .B(\AuI._0637_ ),
    .X(\AuI._0667_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1482_  (.A(\AuI._0664_ ),
    .B(\AuI._0666_ ),
    .C_N(\AuI._0667_ ),
    .X(\AuI._0668_ ));
 sky130_fd_sc_hd__a311o_1 \AuI._1483_  (.A1(\AuI._0645_ ),
    .A2(\AuI._0651_ ),
    .A3(\AuI._0663_ ),
    .B1(\AuI._0668_ ),
    .C1(\AuI._0634_ ),
    .X(\AuI._0669_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1484_  (.A(\AuI._0524_ ),
    .B(\AuI._0527_ ),
    .X(\AuI._0670_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1485_  (.A(\AuI._0524_ ),
    .B(\AuI._0527_ ),
    .Y(\AuI._0671_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1486_  (.A(\AuI._0670_ ),
    .B(\AuI._0671_ ),
    .X(\AuI._0672_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1487_  (.A1(\AuI._0629_ ),
    .A2(\AuI._0644_ ),
    .A3(\AuI._0669_ ),
    .B1(\AuI._0672_ ),
    .X(\AuI._0673_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1488_  (.A(\AuI._0537_ ),
    .B(\AuI._0542_ ),
    .X(\AuI._0674_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1489_  (.A(\AuI._0674_ ),
    .B(\AuI._0670_ ),
    .Y(\AuI._0675_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1490_  (.A(\AuI._0537_ ),
    .B(\AuI._0542_ ),
    .Y(\AuI._0676_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1491_  (.A1(\AuI._0673_ ),
    .A2(\AuI._0675_ ),
    .B1(\AuI._0676_ ),
    .X(\AuI._0677_ ));
 sky130_fd_sc_hd__o221a_1 \AuI._1492_  (.A1(\AuI._0613_ ),
    .A2(\AuI._0614_ ),
    .B1(\AuI._0620_ ),
    .B2(\AuI._0677_ ),
    .C1(\AuI._0615_ ),
    .X(\AuI._0678_ ));
 sky130_fd_sc_hd__or3b_1 \AuI._1493_  (.A(\AuI._0375_ ),
    .B(\AuI._0498_ ),
    .C_N(\AuI._0577_ ),
    .X(\AuI._0679_ ));
 sky130_fd_sc_hd__o21bai_1 \AuI._1494_  (.A1(\AuI._0375_ ),
    .A2(\AuI._0498_ ),
    .B1_N(\AuI._0577_ ),
    .Y(\AuI._0680_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1495_  (.A(\AuI._0679_ ),
    .B(\AuI._0680_ ),
    .Y(\AuI._0681_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1496_  (.A(\AuI._0564_ ),
    .B(\AuI._0566_ ),
    .X(\AuI._0682_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1497_  (.A(\AuI._0564_ ),
    .B(\AuI._0566_ ),
    .Y(\AuI._0683_ ));
 sky130_fd_sc_hd__or2_2 \AuI._1498_  (.A(\AuI._0682_ ),
    .B(\AuI._0683_ ),
    .X(\AuI._0684_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1499_  (.A(\AuI._0680_ ),
    .B(\AuI._0682_ ),
    .Y(\AuI._0685_ ));
 sky130_fd_sc_hd__o311ai_4 \AuI._1500_  (.A1(\AuI._0678_ ),
    .A2(\AuI._0681_ ),
    .A3(\AuI._0684_ ),
    .B1(\AuI._0685_ ),
    .C1(\AuI._0679_ ),
    .Y(\AuI._0686_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1501_  (.A(\AuI._0596_ ),
    .B(\AuI._0598_ ),
    .X(\AuI._0687_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1502_  (.A(\AuI._0583_ ),
    .B(\AuI._0586_ ),
    .X(\AuI._0688_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1503_  (.A(\AuI._0583_ ),
    .B(\AuI._0586_ ),
    .Y(\AuI._0689_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1504_  (.A(\AuI._0688_ ),
    .B(\AuI._0689_ ),
    .Y(\AuI._0690_ ));
 sky130_fd_sc_hd__a21bo_1 \AuI._1505_  (.A1(\AuI._0596_ ),
    .A2(\AuI._0688_ ),
    .B1_N(\AuI._0598_ ),
    .X(\AuI._0691_ ));
 sky130_fd_sc_hd__a31o_2 \AuI._1506_  (.A1(\AuI._0686_ ),
    .A2(\AuI._0687_ ),
    .A3(\AuI._0690_ ),
    .B1(\AuI._0691_ ),
    .X(\AuI._0692_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1507_  (.A(\AuI._0692_ ),
    .X(\AuI._0693_ ));
 sky130_fd_sc_hd__mux2_1 \AuI._1508_  (.A0(\AuI._0608_ ),
    .A1(\AuI._0612_ ),
    .S(\AuI._0693_ ),
    .X(\AuI._0694_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1509_  (.A(\AuI._0599_ ),
    .X(\AuI._0695_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1510_  (.A(\AuI.pe.Significand[0] ),
    .B(\AuI._0695_ ),
    .X(\AuI._0696_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._1511_  (.A(\AuI.operand_a[28] ),
    .B(\AuI.operand_a[29] ),
    .C(\AuI._0604_ ),
    .Y(\AuI._0697_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1512_  (.A(\AuI._0116_ ),
    .B(\AuI._0697_ ),
    .X(\AuI._0698_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1513_  (.A(\AuI._0698_ ),
    .X(\AuI._0699_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1514_  (.A(\AuI._0699_ ),
    .X(\AuI._0700_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1515_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0694_ ),
    .B1(\AuI._0696_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[0] ));
 sky130_fd_sc_hd__buf_2 \AuI._1516_  (.A(\AuI._0692_ ),
    .X(\AuI._0701_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1517_  (.A(\AuI._0599_ ),
    .B(\AuI._0692_ ),
    .Y(\AuI._0702_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1518_  (.A(\AuI._0702_ ),
    .X(\AuI._0703_ ));
 sky130_fd_sc_hd__or2b_1 \AuI._1519_  (.A(\AuI._0656_ ),
    .B_N(\AuI._0653_ ),
    .X(\AuI._0704_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1520_  (.A(\AuI._0704_ ),
    .B(\AuI._0654_ ),
    .Y(\AuI._0705_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1521_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0612_ ),
    .B1(\AuI._0703_ ),
    .B2(\AuI._0705_ ),
    .X(\AuI._0706_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1522_  (.A(\AuI.pe.Significand[1] ),
    .B(\AuI._0695_ ),
    .X(\AuI._0707_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1523_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0706_ ),
    .B1(\AuI._0707_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[1] ));
 sky130_fd_sc_hd__or2_1 \AuI._1524_  (.A(\AuI._0257_ ),
    .B(\AuI._0692_ ),
    .X(\AuI._0708_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1525_  (.A(\AuI._0599_ ),
    .B(\AuI._0692_ ),
    .X(\AuI._0709_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1526_  (.A(\AuI._0709_ ),
    .X(\AuI._0710_ ));
 sky130_fd_sc_hd__a21o_1 \AuI._1527_  (.A1(\AuI._0653_ ),
    .A2(\AuI._0654_ ),
    .B1(\AuI._0656_ ),
    .X(\AuI._0711_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1528_  (.A_N(\AuI._0655_ ),
    .B(\AuI._0652_ ),
    .X(\AuI._0712_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1529_  (.A(\AuI._0711_ ),
    .B(\AuI._0712_ ),
    .Y(\AuI._0713_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1530_  (.A(\AuI._0710_ ),
    .B(\AuI._0713_ ),
    .Y(\AuI._0714_ ));
 sky130_fd_sc_hd__o21ba_1 \AuI._1531_  (.A1(\AuI.pe.Significand[2] ),
    .A2(\AuI._0695_ ),
    .B1_N(\AuI.Exception ),
    .X(\AuI._0715_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1532_  (.A1(\AuI._0708_ ),
    .A2(\AuI._0705_ ),
    .B1(\AuI._0714_ ),
    .C1(\AuI._0715_ ),
    .X(\AuI.result[2] ));
 sky130_fd_sc_hd__inv_2 \AuI._1533_  (.A(\AuI._0713_ ),
    .Y(\AuI._0716_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1534_  (.A(\AuI._0652_ ),
    .B(\AuI._0657_ ),
    .X(\AuI._0717_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1535_  (.A(\AuI._0717_ ),
    .B(\AuI._0658_ ),
    .X(\AuI._0718_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1536_  (.A(\AuI._0702_ ),
    .X(\AuI._0719_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1537_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0716_ ),
    .B1(\AuI._0718_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0720_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1538_  (.A(\AuI._0599_ ),
    .X(\AuI._0721_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1539_  (.A(\AuI.pe.Significand[3] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0722_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1540_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0720_ ),
    .B1(\AuI._0722_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[3] ));
 sky130_fd_sc_hd__a31o_1 \AuI._1541_  (.A1(\AuI._0652_ ),
    .A2(\AuI._0657_ ),
    .A3(\AuI._0658_ ),
    .B1(\AuI._0647_ ),
    .X(\AuI._0723_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1542_  (.A(\AuI._0723_ ),
    .B(\AuI._0659_ ),
    .X(\AuI._0724_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1543_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0718_ ),
    .B1(\AuI._0724_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0725_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1544_  (.A(\AuI.pe.Significand[4] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0726_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1545_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0725_ ),
    .B1(\AuI._0726_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[4] ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1546_  (.A1(\AuI._0649_ ),
    .A2(\AuI._0723_ ),
    .B1(\AuI._0646_ ),
    .Y(\AuI._0727_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1547_  (.A(\AuI._0650_ ),
    .B(\AuI._0727_ ),
    .Y(\AuI._0728_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1548_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0724_ ),
    .B1(\AuI._0728_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0729_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1549_  (.A(\AuI.pe.Significand[5] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0730_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1550_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0729_ ),
    .B1(\AuI._0730_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[5] ));
 sky130_fd_sc_hd__and2b_1 \AuI._1551_  (.A_N(\AuI._0727_ ),
    .B(\AuI._0650_ ),
    .X(\AuI._0731_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1552_  (.A(\AuI._0661_ ),
    .B(\AuI._0731_ ),
    .Y(\AuI._0732_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1553_  (.A(\AuI._0732_ ),
    .B(\AuI._0648_ ),
    .Y(\AuI._0733_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1554_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0728_ ),
    .B1(\AuI._0733_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0734_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1555_  (.A(\AuI.pe.Significand[6] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0735_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1556_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0734_ ),
    .B1(\AuI._0735_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[6] ));
 sky130_fd_sc_hd__a31oi_2 \AuI._1557_  (.A1(\AuI._0645_ ),
    .A2(\AuI._0651_ ),
    .A3(\AuI._0663_ ),
    .B1(\AuI._0666_ ),
    .Y(\AuI._0736_ ));
 sky130_fd_sc_hd__and4_1 \AuI._1558_  (.A(\AuI._0645_ ),
    .B(\AuI._0651_ ),
    .C(\AuI._0663_ ),
    .D(\AuI._0666_ ),
    .X(\AuI._0737_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1559_  (.A(\AuI._0736_ ),
    .B(\AuI._0737_ ),
    .Y(\AuI._0738_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1560_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0733_ ),
    .B1(\AuI._0738_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0739_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1561_  (.A(\AuI.pe.Significand[7] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0740_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1562_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0739_ ),
    .B1(\AuI._0740_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[7] ));
 sky130_fd_sc_hd__nor2_1 \AuI._1563_  (.A(\AuI._0636_ ),
    .B(\AuI._0736_ ),
    .Y(\AuI._0741_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1564_  (.A(\AuI._0667_ ),
    .B(\AuI._0741_ ),
    .Y(\AuI._0742_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1565_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0738_ ),
    .B1(\AuI._0742_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0743_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1566_  (.A(\AuI.pe.Significand[8] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0744_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1567_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0743_ ),
    .B1(\AuI._0744_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[8] ));
 sky130_fd_sc_hd__o31a_1 \AuI._1568_  (.A1(\AuI._0635_ ),
    .A2(\AuI._0636_ ),
    .A3(\AuI._0736_ ),
    .B1(\AuI._0637_ ),
    .X(\AuI._0745_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1569_  (.A(\AuI._0639_ ),
    .B(\AuI._0745_ ),
    .X(\AuI._0746_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1570_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0742_ ),
    .B1(\AuI._0746_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0747_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1571_  (.A(\AuI.pe.Significand[9] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0748_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1572_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0747_ ),
    .B1(\AuI._0748_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[9] ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1573_  (.A1(\AuI._0639_ ),
    .A2(\AuI._0745_ ),
    .B1(\AuI._0641_ ),
    .Y(\AuI._0749_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1574_  (.A(\AuI._0638_ ),
    .B(\AuI._0749_ ),
    .Y(\AuI._0750_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1575_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0746_ ),
    .B1(\AuI._0750_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0751_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1576_  (.A(\AuI.pe.Significand[10] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0752_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1577_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0751_ ),
    .B1(\AuI._0752_ ),
    .C1(\AuI._0700_ ),
    .X(\AuI.result[10] ));
 sky130_fd_sc_hd__and3_1 \AuI._1578_  (.A(\AuI._0638_ ),
    .B(\AuI._0639_ ),
    .C(\AuI._0667_ ),
    .X(\AuI._0753_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1579_  (.A1(\AuI._0736_ ),
    .A2(\AuI._0753_ ),
    .B1(\AuI._0643_ ),
    .Y(\AuI._0754_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1580_  (.A_N(\AuI._0754_ ),
    .B(\AuI._0633_ ),
    .X(\AuI._0755_ ));
 sky130_fd_sc_hd__and2b_1 \AuI._1581_  (.A_N(\AuI._0633_ ),
    .B(\AuI._0754_ ),
    .X(\AuI._0756_ ));
 sky130_fd_sc_hd__nor2_1 \AuI._1582_  (.A(\AuI._0755_ ),
    .B(\AuI._0756_ ),
    .Y(\AuI._0757_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1583_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0750_ ),
    .B1(\AuI._0757_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0758_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1584_  (.A(\AuI.pe.Significand[11] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0759_ ));
 sky130_fd_sc_hd__buf_2 \AuI._1585_  (.A(\AuI._0699_ ),
    .X(\AuI._0760_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1586_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0758_ ),
    .B1(\AuI._0759_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[11] ));
 sky130_fd_sc_hd__or2_1 \AuI._1587_  (.A(\AuI._0630_ ),
    .B(\AuI._0623_ ),
    .X(\AuI._0761_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1588_  (.A(\AuI._0624_ ),
    .B(\AuI._0755_ ),
    .X(\AuI._0762_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1589_  (.A(\AuI._0761_ ),
    .B(\AuI._0762_ ),
    .Y(\AuI._0763_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1590_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0757_ ),
    .B1(\AuI._0763_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0764_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1591_  (.A(\AuI.pe.Significand[12] ),
    .B(\AuI._0721_ ),
    .X(\AuI._0765_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1592_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0764_ ),
    .B1(\AuI._0765_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[12] ));
 sky130_fd_sc_hd__o31a_1 \AuI._1593_  (.A1(\AuI._0623_ ),
    .A2(\AuI._0624_ ),
    .A3(\AuI._0755_ ),
    .B1(\AuI._0627_ ),
    .X(\AuI._0766_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1594_  (.A(\AuI._0626_ ),
    .B(\AuI._0766_ ),
    .X(\AuI._0767_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1595_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0763_ ),
    .B1(\AuI._0767_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0768_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI._1596_  (.A(\AuI._0599_ ),
    .X(\AuI._0769_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1597_  (.A(\AuI.pe.Significand[13] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0770_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1598_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0768_ ),
    .B1(\AuI._0770_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[13] ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1599_  (.A1(\AuI._0626_ ),
    .A2(\AuI._0766_ ),
    .B1(\AuI._0621_ ),
    .Y(\AuI._0771_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1600_  (.A(\AuI._0625_ ),
    .B(\AuI._0771_ ),
    .Y(\AuI._0772_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1601_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0767_ ),
    .B1(\AuI._0772_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0773_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1602_  (.A(\AuI.pe.Significand[14] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0774_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1603_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0773_ ),
    .B1(\AuI._0774_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[14] ));
 sky130_fd_sc_hd__nand4_1 \AuI._1604_  (.A(\AuI._0629_ ),
    .B(\AuI._0644_ ),
    .C(\AuI._0669_ ),
    .D(\AuI._0672_ ),
    .Y(\AuI._0775_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1605_  (.A(\AuI._0673_ ),
    .B(\AuI._0775_ ),
    .Y(\AuI._0776_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1606_  (.A(\AuI._0710_ ),
    .B(\AuI._0776_ ),
    .Y(\AuI._0777_ ));
 sky130_fd_sc_hd__o21ba_1 \AuI._1607_  (.A1(\AuI.pe.Significand[15] ),
    .A2(\AuI._0695_ ),
    .B1_N(\AuI.Exception ),
    .X(\AuI._0778_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1608_  (.A1(\AuI._0708_ ),
    .A2(\AuI._0772_ ),
    .B1(\AuI._0777_ ),
    .C1(\AuI._0778_ ),
    .X(\AuI.result[15] ));
 sky130_fd_sc_hd__or2b_1 \AuI._1609_  (.A(\AuI._0670_ ),
    .B_N(\AuI._0673_ ),
    .X(\AuI._0779_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1610_  (.A(\AuI._0676_ ),
    .B(\AuI._0674_ ),
    .X(\AuI._0780_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1611_  (.A(\AuI._0779_ ),
    .B(\AuI._0780_ ),
    .Y(\AuI._0781_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1612_  (.A(\AuI._0769_ ),
    .B(\AuI._0776_ ),
    .Y(\AuI._0782_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._1613_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0781_ ),
    .B1(\AuI._0782_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0783_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1614_  (.A1(\AuI.pe.Significand[16] ),
    .A2(\AuI._0695_ ),
    .B1(\AuI._0760_ ),
    .C1(\AuI._0783_ ),
    .X(\AuI.result[16] ));
 sky130_fd_sc_hd__xor2_1 \AuI._1615_  (.A(\AuI._0677_ ),
    .B(\AuI._0619_ ),
    .X(\AuI._0784_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1616_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0781_ ),
    .B1(\AuI._0784_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0785_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1617_  (.A(\AuI.pe.Significand[17] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0786_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1618_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0785_ ),
    .B1(\AuI._0786_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[17] ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1619_  (.A1(\AuI._0677_ ),
    .A2(\AuI._0619_ ),
    .B1(\AuI._0614_ ),
    .Y(\AuI._0787_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI._1620_  (.A(\AuI._0617_ ),
    .B(\AuI._0787_ ),
    .Y(\AuI._0788_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1621_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0784_ ),
    .B1(\AuI._0788_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0789_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1622_  (.A(\AuI.pe.Significand[18] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0790_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1623_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0789_ ),
    .B1(\AuI._0790_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[18] ));
 sky130_fd_sc_hd__xor2_1 \AuI._1624_  (.A(\AuI._0678_ ),
    .B(\AuI._0684_ ),
    .X(\AuI._0791_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1625_  (.A(\AuI._0258_ ),
    .B(\AuI._0788_ ),
    .X(\AuI._0792_ ));
 sky130_fd_sc_hd__a22o_1 \AuI._1626_  (.A1(\AuI._0701_ ),
    .A2(\AuI._0791_ ),
    .B1(\AuI._0792_ ),
    .B2(\AuI._0719_ ),
    .X(\AuI._0793_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1627_  (.A1(\AuI.pe.Significand[19] ),
    .A2(\AuI._0695_ ),
    .B1(\AuI._0760_ ),
    .C1(\AuI._0793_ ),
    .X(\AuI.result[19] ));
 sky130_fd_sc_hd__o21ba_1 \AuI._1628_  (.A1(\AuI._0678_ ),
    .A2(\AuI._0684_ ),
    .B1_N(\AuI._0682_ ),
    .X(\AuI._0794_ ));
 sky130_fd_sc_hd__xor2_1 \AuI._1629_  (.A(\AuI._0681_ ),
    .B(\AuI._0794_ ),
    .X(\AuI._0795_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1630_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0791_ ),
    .B1(\AuI._0795_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0796_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1631_  (.A(\AuI.pe.Significand[20] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0797_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1632_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0796_ ),
    .B1(\AuI._0797_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[20] ));
 sky130_fd_sc_hd__xor2_1 \AuI._1633_  (.A(\AuI._0686_ ),
    .B(\AuI._0690_ ),
    .X(\AuI._0798_ ));
 sky130_fd_sc_hd__o22a_1 \AuI._1634_  (.A1(\AuI._0693_ ),
    .A2(\AuI._0795_ ),
    .B1(\AuI._0798_ ),
    .B2(\AuI._0703_ ),
    .X(\AuI._0799_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1635_  (.A(\AuI.pe.Significand[21] ),
    .B(\AuI._0769_ ),
    .X(\AuI._0800_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1636_  (.A1(\AuI._0259_ ),
    .A2(\AuI._0799_ ),
    .B1(\AuI._0800_ ),
    .C1(\AuI._0760_ ),
    .X(\AuI.result[21] ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1637_  (.A1(\AuI._0686_ ),
    .A2(\AuI._0690_ ),
    .B1(\AuI._0688_ ),
    .Y(\AuI._0801_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1638_  (.A1(\AuI._0687_ ),
    .A2(\AuI._0801_ ),
    .B1(\AuI._0710_ ),
    .Y(\AuI._0802_ ));
 sky130_fd_sc_hd__o221a_1 \AuI._1639_  (.A1(\AuI.pe.Significand[22] ),
    .A2(\AuI._0599_ ),
    .B1(\AuI._0708_ ),
    .B2(\AuI._0798_ ),
    .C1(\AuI._0698_ ),
    .X(\AuI._0803_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1640_  (.A(\AuI._0802_ ),
    .B(\AuI._0803_ ),
    .X(\AuI._0804_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI._1641_  (.A(\AuI._0804_ ),
    .X(\AuI.result[22] ));
 sky130_fd_sc_hd__o221a_1 \AuI._1642_  (.A1(\AuI.exponent_sub[0] ),
    .A2(\AuI._0769_ ),
    .B1(\AuI._0708_ ),
    .B2(\AuI.exp_a ),
    .C1(\AuI._0699_ ),
    .X(\AuI._0000_ ));
 sky130_fd_sc_hd__a21boi_1 \AuI._1643_  (.A1(\AuI.exp_a ),
    .A2(\AuI._0710_ ),
    .B1_N(\AuI._0000_ ),
    .Y(\AuI.result[23] ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1644_  (.A1(\AuI.exp_a ),
    .A2(\AuI._0710_ ),
    .B1(\AuI.operand_a[24] ),
    .Y(\AuI._0001_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1645_  (.A1(\AuI.exponent_sub[1] ),
    .A2(\AuI._0769_ ),
    .B1(\AuI._0699_ ),
    .Y(\AuI._0002_ ));
 sky130_fd_sc_hd__a31o_1 \AuI._1646_  (.A1(\AuI.exp_a ),
    .A2(\AuI.operand_a[24] ),
    .A3(\AuI._0710_ ),
    .B1(\AuI._0002_ ),
    .X(\AuI._0003_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI._1647_  (.A1(\AuI._0695_ ),
    .A2(\AuI._0001_ ),
    .B1(\AuI._0003_ ),
    .Y(\AuI.result[24] ));
 sky130_fd_sc_hd__a31o_1 \AuI._1648_  (.A1(\AuI.exp_a ),
    .A2(\AuI.operand_a[24] ),
    .A3(\AuI._0710_ ),
    .B1(\AuI.operand_a[25] ),
    .X(\AuI._0004_ ));
 sky130_fd_sc_hd__o221a_1 \AuI._1649_  (.A1(\AuI.exponent_sub[2] ),
    .A2(\AuI._0695_ ),
    .B1(\AuI._0602_ ),
    .B2(\AuI._0719_ ),
    .C1(\AuI._0699_ ),
    .X(\AuI._0005_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1650_  (.A1(\AuI._0606_ ),
    .A2(\AuI._0004_ ),
    .B1(\AuI._0005_ ),
    .X(\AuI.result[25] ));
 sky130_fd_sc_hd__a211o_1 \AuI._1651_  (.A1(\AuI._0603_ ),
    .A2(\AuI._0692_ ),
    .B1(\AuI.operand_a[26] ),
    .C1(\AuI._0258_ ),
    .X(\AuI._0006_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1652_  (.A1(\AuI.exponent_sub[3] ),
    .A2(\AuI._0769_ ),
    .B1(\AuI._0699_ ),
    .X(\AuI._0007_ ));
 sky130_fd_sc_hd__and2_1 \AuI._1653_  (.A(\AuI.operand_a[26] ),
    .B(\AuI._0603_ ),
    .X(\AuI._0008_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1654_  (.A(\AuI._0008_ ),
    .B(\AuI._0710_ ),
    .Y(\AuI._0009_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1655_  (.A(\AuI._0006_ ),
    .B(\AuI._0007_ ),
    .C(\AuI._0009_ ),
    .X(\AuI._0010_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI._1656_  (.A(\AuI._0010_ ),
    .X(\AuI.result[26] ));
 sky130_fd_sc_hd__a211o_1 \AuI._1657_  (.A1(\AuI._0008_ ),
    .A2(\AuI._0692_ ),
    .B1(\AuI.operand_a[27] ),
    .C1(\AuI._0258_ ),
    .X(\AuI._0011_ ));
 sky130_fd_sc_hd__nand2_1 \AuI._1658_  (.A(\AuI._0604_ ),
    .B(\AuI._0710_ ),
    .Y(\AuI._0012_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1659_  (.A1(\AuI.exponent_sub[4] ),
    .A2(\AuI._0599_ ),
    .B1(\AuI._0698_ ),
    .X(\AuI._0013_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1660_  (.A(\AuI._0011_ ),
    .B(\AuI._0012_ ),
    .C(\AuI._0013_ ),
    .X(\AuI._0014_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI._1661_  (.A(\AuI._0014_ ),
    .X(\AuI.result[27] ));
 sky130_fd_sc_hd__a211o_1 \AuI._1662_  (.A1(\AuI._0604_ ),
    .A2(\AuI._0692_ ),
    .B1(\AuI.operand_a[28] ),
    .C1(\AuI._0258_ ),
    .X(\AuI._0015_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1663_  (.A1(\AuI.exponent_sub[5] ),
    .A2(\AuI._0599_ ),
    .B1(\AuI._0699_ ),
    .X(\AuI._0016_ ));
 sky130_fd_sc_hd__nand3_1 \AuI._1664_  (.A(\AuI.operand_a[28] ),
    .B(\AuI._0604_ ),
    .C(\AuI._0710_ ),
    .Y(\AuI._0017_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1665_  (.A(\AuI._0015_ ),
    .B(\AuI._0016_ ),
    .C(\AuI._0017_ ),
    .X(\AuI._0018_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI._1666_  (.A(\AuI._0018_ ),
    .X(\AuI.result[28] ));
 sky130_fd_sc_hd__a311o_1 \AuI._1667_  (.A1(\AuI.operand_a[28] ),
    .A2(\AuI._0604_ ),
    .A3(\AuI._0692_ ),
    .B1(\AuI.operand_a[29] ),
    .C1(\AuI._0258_ ),
    .X(\AuI._0019_ ));
 sky130_fd_sc_hd__o21a_1 \AuI._1668_  (.A1(\AuI.exponent_sub[6] ),
    .A2(\AuI._0599_ ),
    .B1(\AuI._0699_ ),
    .X(\AuI._0020_ ));
 sky130_fd_sc_hd__or2_1 \AuI._1669_  (.A(\AuI._0702_ ),
    .B(\AuI._0697_ ),
    .X(\AuI._0021_ ));
 sky130_fd_sc_hd__and3_1 \AuI._1670_  (.A(\AuI._0019_ ),
    .B(\AuI._0020_ ),
    .C(\AuI._0021_ ),
    .X(\AuI._0022_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI._1671_  (.A(\AuI._0022_ ),
    .X(\AuI.result[29] ));
 sky130_fd_sc_hd__o21ai_1 \AuI._1672_  (.A1(\AuI.exponent_sub[7] ),
    .A2(\AuI._0695_ ),
    .B1(\AuI._0699_ ),
    .Y(\AuI._0023_ ));
 sky130_fd_sc_hd__a31oi_1 \AuI._1673_  (.A1(\AuI._0116_ ),
    .A2(\AuI._0695_ ),
    .A3(\AuI._0021_ ),
    .B1(\AuI._0023_ ),
    .Y(\AuI.result[30] ));
 sky130_fd_sc_hd__or3_1 \AuI._1674_  (.A(\AuI._0119_ ),
    .B(\AuI._0120_ ),
    .C(\AuI._0138_ ),
    .X(\AuI._0024_ ));
 sky130_fd_sc_hd__o211a_1 \AuI._1675_  (.A1(net29),
    .A2(\AuI._0126_ ),
    .B1(\AuI._0699_ ),
    .C1(\AuI._0024_ ),
    .X(\AuI.result[31] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._400_  (.A(\AuI.pe.significand[16] ),
    .X(\AuI.pe._367_ ));
 sky130_fd_sc_hd__or4b_4 \AuI.pe._401_  (.A(\AuI.pe.significand[21] ),
    .B(\AuI.pe.significand[23] ),
    .C(\AuI.pe.significand[22] ),
    .D_N(\AuI.pe.significand[24] ),
    .X(\AuI.pe._368_ ));
 sky130_fd_sc_hd__or4_2 \AuI.pe._402_  (.A(\AuI.pe.significand[17] ),
    .B(\AuI.pe.significand[18] ),
    .C(\AuI.pe.significand[19] ),
    .D(\AuI.pe.significand[20] ),
    .X(\AuI.pe._369_ ));
 sky130_fd_sc_hd__or3_4 \AuI.pe._403_  (.A(\AuI.pe._367_ ),
    .B(\AuI.pe._368_ ),
    .C(\AuI.pe._369_ ),
    .X(\AuI.pe._370_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._404_  (.A(\AuI.pe.significand[12] ),
    .B(\AuI.pe.significand[13] ),
    .C(\AuI.pe.significand[14] ),
    .D(\AuI.pe.significand[15] ),
    .X(\AuI.pe._371_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._405_  (.A(\AuI.pe._371_ ),
    .X(\AuI.pe._372_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._406_  (.A(\AuI.pe.significand[9] ),
    .B(\AuI.pe.significand[10] ),
    .C(\AuI.pe.significand[11] ),
    .X(\AuI.pe._373_ ));
 sky130_fd_sc_hd__or3_2 \AuI.pe._407_  (.A(\AuI.pe.significand[8] ),
    .B(\AuI.pe._372_ ),
    .C(\AuI.pe._373_ ),
    .X(\AuI.pe._374_ ));
 sky130_fd_sc_hd__or4_2 \AuI.pe._408_  (.A(\AuI.pe.significand[5] ),
    .B(\AuI.pe.significand[4] ),
    .C(\AuI.pe.significand[6] ),
    .D(\AuI.pe.significand[7] ),
    .X(\AuI.pe._375_ ));
 sky130_fd_sc_hd__or2b_1 \AuI.pe._409_  (.A(\AuI.pe.significand[3] ),
    .B_N(\AuI.pe.significand[2] ),
    .X(\AuI.pe._376_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._410_  (.A(\AuI.pe._370_ ),
    .B(\AuI.pe._374_ ),
    .C(\AuI.pe._375_ ),
    .D(\AuI.pe._376_ ),
    .X(\AuI.pe._377_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._411_  (.A(\AuI.pe.significand[11] ),
    .X(\AuI.pe._378_ ));
 sky130_fd_sc_hd__or4_2 \AuI.pe._412_  (.A(\AuI.pe._367_ ),
    .B(\AuI.pe._368_ ),
    .C(\AuI.pe._369_ ),
    .D(\AuI.pe._372_ ),
    .X(\AuI.pe._379_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._413_  (.A(\AuI.pe.significand[10] ),
    .X(\AuI.pe._380_ ));
 sky130_fd_sc_hd__or3b_1 \AuI.pe._414_  (.A(\AuI.pe._378_ ),
    .B(\AuI.pe._379_ ),
    .C_N(\AuI.pe._380_ ),
    .X(\AuI.pe._381_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._415_  (.A(\AuI.pe.significand[16] ),
    .Y(\AuI.pe._382_ ));
 sky130_fd_sc_hd__nor4b_1 \AuI.pe._416_  (.A(\AuI.pe.significand[21] ),
    .B(\AuI.pe.significand[23] ),
    .C(\AuI.pe.significand[22] ),
    .D_N(\AuI.pe.significand[24] ),
    .Y(\AuI.pe._383_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI.pe._417_  (.A(\AuI.pe._383_ ),
    .X(\AuI.pe._384_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._418_  (.A(\AuI.pe.significand[18] ),
    .X(\AuI.pe._385_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._419_  (.A(\AuI.pe.significand[19] ),
    .X(\AuI.pe._386_ ));
 sky130_fd_sc_hd__nor4_4 \AuI.pe._420_  (.A(\AuI.pe.significand[17] ),
    .B(\AuI.pe._385_ ),
    .C(\AuI.pe._386_ ),
    .D(\AuI.pe.significand[20] ),
    .Y(\AuI.pe._387_ ));
 sky130_fd_sc_hd__and3_2 \AuI.pe._421_  (.A(\AuI.pe._382_ ),
    .B(\AuI.pe._384_ ),
    .C(\AuI.pe._387_ ),
    .X(\AuI.pe._388_ ));
 sky130_fd_sc_hd__nor3_1 \AuI.pe._422_  (.A(\AuI.pe.significand[13] ),
    .B(\AuI.pe.significand[14] ),
    .C(\AuI.pe.significand[15] ),
    .Y(\AuI.pe._389_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._423_  (.A_N(\AuI.pe.significand[15] ),
    .B(\AuI.pe.significand[14] ),
    .X(\AuI.pe._390_ ));
 sky130_fd_sc_hd__and4_2 \AuI.pe._424_  (.A(\AuI.pe._382_ ),
    .B(\AuI.pe._384_ ),
    .C(\AuI.pe._387_ ),
    .D(\AuI.pe._390_ ),
    .X(\AuI.pe._391_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._425_  (.A1(\AuI.pe.significand[12] ),
    .A2(\AuI.pe._388_ ),
    .A3(\AuI.pe._389_ ),
    .B1(\AuI.pe._391_ ),
    .X(\AuI.pe._392_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._426_  (.A(\AuI.pe.significand[8] ),
    .X(\AuI.pe._393_ ));
 sky130_fd_sc_hd__nor3_1 \AuI.pe._427_  (.A(\AuI.pe.significand[9] ),
    .B(\AuI.pe.significand[10] ),
    .C(\AuI.pe.significand[11] ),
    .Y(\AuI.pe._394_ ));
 sky130_fd_sc_hd__nor4_4 \AuI.pe._428_  (.A(\AuI.pe._367_ ),
    .B(\AuI.pe._368_ ),
    .C(\AuI.pe._369_ ),
    .D(\AuI.pe._372_ ),
    .Y(\AuI.pe._395_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._429_  (.A(\AuI.pe._393_ ),
    .B(\AuI.pe._394_ ),
    .C(\AuI.pe._395_ ),
    .X(\AuI.pe._396_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._430_  (.A(\AuI.pe._396_ ),
    .X(\AuI.pe._397_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._431_  (.A(\AuI.pe._392_ ),
    .B(\AuI.pe._397_ ),
    .Y(\AuI.pe._398_ ));
 sky130_fd_sc_hd__and3_2 \AuI.pe._432_  (.A(\AuI.pe._367_ ),
    .B(\AuI.pe._384_ ),
    .C(\AuI.pe._387_ ),
    .X(\AuI.pe._399_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._433_  (.A(\AuI.pe.significand[20] ),
    .Y(\AuI.pe._000_ ));
 sky130_fd_sc_hd__and4b_1 \AuI.pe._434_  (.A_N(\AuI.pe._386_ ),
    .B(\AuI.pe._000_ ),
    .C(\AuI.pe._383_ ),
    .D(\AuI.pe._385_ ),
    .X(\AuI.pe._001_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._435_  (.A(\AuI.pe._001_ ),
    .X(\AuI.pe._002_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._436_  (.A(\AuI.pe._000_ ),
    .B(\AuI.pe._368_ ),
    .Y(\AuI.pe._003_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._437_  (.A(\AuI.pe._003_ ),
    .X(\AuI.pe._004_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._438_  (.A_N(\AuI.pe.significand[23] ),
    .B(\AuI.pe.significand[24] ),
    .X(\AuI.pe._005_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._439_  (.A(\AuI.pe.significand[22] ),
    .B(\AuI.pe._005_ ),
    .X(\AuI.pe._006_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._440_  (.A(\AuI.pe._399_ ),
    .B(\AuI.pe._002_ ),
    .C(\AuI.pe._004_ ),
    .D(\AuI.pe._006_ ),
    .X(\AuI.pe._007_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._441_  (.A(\AuI.pe.significand[8] ),
    .Y(\AuI.pe._008_ ));
 sky130_fd_sc_hd__and3b_1 \AuI.pe._442_  (.A_N(\AuI.pe._372_ ),
    .B(\AuI.pe._394_ ),
    .C(\AuI.pe._008_ ),
    .X(\AuI.pe._009_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._443_  (.A(\AuI.pe.significand[6] ),
    .B(\AuI.pe.significand[7] ),
    .Y(\AuI.pe._010_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._444_  (.A_N(\AuI.pe.significand[5] ),
    .B(\AuI.pe._010_ ),
    .X(\AuI.pe._011_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._445_  (.A(\AuI.pe.significand[4] ),
    .B(\AuI.pe._388_ ),
    .C(\AuI.pe._009_ ),
    .D(\AuI.pe._011_ ),
    .X(\AuI.pe._012_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._446_  (.A(\AuI.pe.significand[1] ),
    .X(\AuI.pe._013_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._447_  (.A(\AuI.pe.significand[0] ),
    .X(\AuI.pe._014_ ));
 sky130_fd_sc_hd__or4b_1 \AuI.pe._448_  (.A(\AuI.pe._013_ ),
    .B(\AuI.pe.significand[2] ),
    .C(\AuI.pe.significand[3] ),
    .D_N(\AuI.pe._014_ ),
    .X(\AuI.pe._015_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._449_  (.A(\AuI.pe._370_ ),
    .B(\AuI.pe._374_ ),
    .C(\AuI.pe._375_ ),
    .D(\AuI.pe._015_ ),
    .X(\AuI.pe._016_ ));
 sky130_fd_sc_hd__or4b_1 \AuI.pe._450_  (.A(\AuI.pe.significand[7] ),
    .B(\AuI.pe._370_ ),
    .C(\AuI.pe._374_ ),
    .D_N(\AuI.pe.significand[6] ),
    .X(\AuI.pe._017_ ));
 sky130_fd_sc_hd__and4bb_1 \AuI.pe._451_  (.A_N(\AuI.pe._007_ ),
    .B_N(\AuI.pe._012_ ),
    .C(\AuI.pe._016_ ),
    .D(\AuI.pe._017_ ),
    .X(\AuI.pe._018_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._452_  (.A(\AuI.pe._377_ ),
    .B(\AuI.pe._381_ ),
    .C(\AuI.pe._398_ ),
    .D(\AuI.pe._018_ ),
    .X(\AuI.pe._019_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._453_  (.A(\AuI.exp_a ),
    .B(\AuI.pe._019_ ),
    .Y(\AuI.exponent_sub[0] ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._454_  (.A(\AuI.pe._014_ ),
    .X(\AuI.pe._020_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._455_  (.A_N(\AuI.pe._005_ ),
    .B(\AuI.pe._020_ ),
    .X(\AuI.pe._021_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI.pe._456_  (.A(\AuI.pe._021_ ),
    .X(\AuI.pe.Significand[0] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._457_  (.A(\AuI.pe._006_ ),
    .X(\AuI.pe._022_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._458_  (.A(\AuI.pe._022_ ),
    .X(\AuI.pe._023_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._459_  (.A(\AuI.pe.significand[24] ),
    .X(\AuI.pe._024_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._460_  (.A(\AuI.pe.significand[23] ),
    .X(\AuI.pe._025_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._461_  (.A(\AuI.pe._025_ ),
    .X(\AuI.pe._026_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._462_  (.A(\AuI.pe._024_ ),
    .B(\AuI.pe._026_ ),
    .X(\AuI.pe._027_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._463_  (.A(\AuI.pe._013_ ),
    .X(\AuI.pe._028_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._464_  (.A(\AuI.pe._028_ ),
    .X(\AuI.pe._029_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._465_  (.A(\AuI.pe._014_ ),
    .X(\AuI.pe._030_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._466_  (.A1(\AuI.pe._028_ ),
    .A2(\AuI.pe._030_ ),
    .B1(\AuI.pe._024_ ),
    .Y(\AuI.pe._031_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._467_  (.A1(\AuI.pe._029_ ),
    .A2(\AuI.pe._020_ ),
    .B1(\AuI.pe._031_ ),
    .X(\AuI.pe._032_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._468_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._027_ ),
    .B2(\AuI.pe._029_ ),
    .C1(\AuI.pe._032_ ),
    .X(\AuI.pe.Significand[1] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._469_  (.A(\AuI.pe.significand[2] ),
    .X(\AuI.pe._033_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._470_  (.A1(\AuI.pe._028_ ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._027_ ),
    .B2(\AuI.pe._033_ ),
    .X(\AuI.pe._034_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._471_  (.A(\AuI.pe.significand[24] ),
    .Y(\AuI.pe._035_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._472_  (.A(\AuI.pe._035_ ),
    .X(\AuI.pe._036_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._473_  (.A(\AuI.pe._036_ ),
    .X(\AuI.pe._037_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._474_  (.A(\AuI.pe._013_ ),
    .B(\AuI.pe._014_ ),
    .C(\AuI.pe.significand[2] ),
    .X(\AuI.pe._038_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._475_  (.A1(\AuI.pe._013_ ),
    .A2(\AuI.pe._014_ ),
    .B1(\AuI.pe._033_ ),
    .Y(\AuI.pe._039_ ));
 sky130_fd_sc_hd__and3b_1 \AuI.pe._476_  (.A_N(\AuI.pe.significand[22] ),
    .B(\AuI.pe._005_ ),
    .C(\AuI.pe.significand[21] ),
    .X(\AuI.pe._040_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._477_  (.A(\AuI.pe._040_ ),
    .X(\AuI.pe._041_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._478_  (.A(\AuI.pe._041_ ),
    .X(\AuI.pe._042_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._479_  (.A1(\AuI.pe._037_ ),
    .A2(\AuI.pe._038_ ),
    .A3(\AuI.pe._039_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._030_ ),
    .X(\AuI.pe._043_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._480_  (.A(\AuI.pe._034_ ),
    .B(\AuI.pe._043_ ),
    .X(\AuI.pe._044_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI.pe._481_  (.A(\AuI.pe._044_ ),
    .X(\AuI.pe.Significand[2] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._482_  (.A(\AuI.pe.significand[3] ),
    .X(\AuI.pe._045_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._483_  (.A(\AuI.pe._045_ ),
    .X(\AuI.pe._046_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._484_  (.A(\AuI.pe._046_ ),
    .B(\AuI.pe._038_ ),
    .Y(\AuI.pe._047_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._485_  (.A(\AuI.pe.significand[1] ),
    .B(\AuI.pe.significand[0] ),
    .C(\AuI.pe.significand[2] ),
    .D(\AuI.pe.significand[3] ),
    .X(\AuI.pe._048_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI.pe._486_  (.A(\AuI.pe._048_ ),
    .X(\AuI.pe._049_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._487_  (.A(\AuI.pe._004_ ),
    .X(\AuI.pe._050_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._488_  (.A1(\AuI.pe._033_ ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._027_ ),
    .B2(\AuI.pe._045_ ),
    .X(\AuI.pe._051_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._489_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._029_ ),
    .C1(\AuI.pe._051_ ),
    .X(\AuI.pe._052_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._490_  (.A1(\AuI.pe._037_ ),
    .A2(\AuI.pe._047_ ),
    .A3(\AuI.pe._049_ ),
    .B1(\AuI.pe._052_ ),
    .X(\AuI.pe.Significand[3] ));
 sky130_fd_sc_hd__and3_2 \AuI.pe._491_  (.A(\AuI.pe._386_ ),
    .B(\AuI.pe._000_ ),
    .C(\AuI.pe._384_ ),
    .X(\AuI.pe._053_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._492_  (.A(\AuI.pe._053_ ),
    .X(\AuI.pe._054_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._493_  (.A(\AuI.pe._033_ ),
    .X(\AuI.pe._055_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._494_  (.A(\AuI.pe.significand[4] ),
    .X(\AuI.pe._056_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._495_  (.A1(\AuI.pe._045_ ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._027_ ),
    .B2(\AuI.pe._056_ ),
    .X(\AuI.pe._057_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._496_  (.A1(\AuI.pe._028_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._055_ ),
    .C1(\AuI.pe._057_ ),
    .X(\AuI.pe._058_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._497_  (.A(\AuI.pe._056_ ),
    .X(\AuI.pe._059_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._498_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._049_ ),
    .B1(\AuI.pe._024_ ),
    .Y(\AuI.pe._060_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._499_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._049_ ),
    .B1(\AuI.pe._060_ ),
    .X(\AuI.pe._061_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._500_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._054_ ),
    .B1(\AuI.pe._058_ ),
    .C1(\AuI.pe._061_ ),
    .X(\AuI.pe.Significand[4] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._501_  (.A(\AuI.pe.significand[5] ),
    .X(\AuI.pe._062_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._502_  (.A(\AuI.pe._062_ ),
    .X(\AuI.pe._063_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._503_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._049_ ),
    .B1(\AuI.pe._063_ ),
    .Y(\AuI.pe._064_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._504_  (.A(\AuI.pe.significand[5] ),
    .B(\AuI.pe.significand[4] ),
    .C(\AuI.pe._049_ ),
    .X(\AuI.pe._065_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._505_  (.A(\AuI.pe._002_ ),
    .X(\AuI.pe._066_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._506_  (.A1(\AuI.pe.significand[4] ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._027_ ),
    .B2(\AuI.pe._062_ ),
    .X(\AuI.pe._067_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._507_  (.A1(\AuI.pe._033_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._045_ ),
    .C1(\AuI.pe._067_ ),
    .X(\AuI.pe._068_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._508_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._029_ ),
    .C1(\AuI.pe._068_ ),
    .X(\AuI.pe._069_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._509_  (.A1(\AuI.pe._037_ ),
    .A2(\AuI.pe._064_ ),
    .A3(\AuI.pe._065_ ),
    .B1(\AuI.pe._069_ ),
    .X(\AuI.pe.Significand[5] ));
 sky130_fd_sc_hd__or2_2 \AuI.pe._510_  (.A(\AuI.pe.significand[6] ),
    .B(\AuI.pe._065_ ),
    .X(\AuI.pe._070_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._511_  (.A(\AuI.pe.significand[6] ),
    .X(\AuI.pe._071_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._512_  (.A(\AuI.pe._071_ ),
    .X(\AuI.pe._072_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._513_  (.A(\AuI.pe._072_ ),
    .B(\AuI.pe._065_ ),
    .Y(\AuI.pe._073_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._514_  (.A(\AuI.pe._024_ ),
    .X(\AuI.pe._074_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._515_  (.A1(\AuI.pe._070_ ),
    .A2(\AuI.pe._073_ ),
    .B1(\AuI.pe._074_ ),
    .Y(\AuI.pe._075_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._516_  (.A(\AuI.pe._385_ ),
    .B(\AuI.pe._386_ ),
    .Y(\AuI.pe._076_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._517_  (.A(\AuI.pe.significand[17] ),
    .B(\AuI.pe._000_ ),
    .C(\AuI.pe._383_ ),
    .D(\AuI.pe._076_ ),
    .X(\AuI.pe._077_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._518_  (.A(\AuI.pe._077_ ),
    .X(\AuI.pe._078_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._519_  (.A(\AuI.pe._078_ ),
    .X(\AuI.pe._079_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._520_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._022_ ),
    .B2(\AuI.pe._062_ ),
    .C1(\AuI.pe._037_ ),
    .X(\AuI.pe._080_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._521_  (.A1(\AuI.pe.significand[3] ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._056_ ),
    .C1(\AuI.pe._080_ ),
    .X(\AuI.pe._081_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._522_  (.A1(\AuI.pe._028_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._055_ ),
    .C1(\AuI.pe._081_ ),
    .X(\AuI.pe._082_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._523_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._079_ ),
    .B1(\AuI.pe._082_ ),
    .Y(\AuI.pe._083_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._524_  (.A(\AuI.pe._075_ ),
    .B(\AuI.pe._083_ ),
    .Y(\AuI.pe.Significand[6] ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._525_  (.A(\AuI.pe.significand[7] ),
    .X(\AuI.pe._084_ ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._526_  (.A(\AuI.pe._084_ ),
    .B(\AuI.pe._070_ ),
    .X(\AuI.pe._085_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._527_  (.A(\AuI.pe._399_ ),
    .X(\AuI.pe._086_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._528_  (.A1(\AuI.pe._014_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._066_ ),
    .B2(\AuI.pe._033_ ),
    .X(\AuI.pe._087_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._529_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._054_ ),
    .B1(\AuI.pe._087_ ),
    .X(\AuI.pe._088_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._530_  (.A(\AuI.pe.significand[7] ),
    .X(\AuI.pe._089_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._531_  (.A1(\AuI.pe._089_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._037_ ),
    .X(\AuI.pe._090_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._532_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._023_ ),
    .B2(\AuI.pe._072_ ),
    .C1(\AuI.pe._090_ ),
    .X(\AuI.pe._091_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._533_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._042_ ),
    .B1(\AuI.pe._079_ ),
    .B2(\AuI.pe._029_ ),
    .C1(\AuI.pe._091_ ),
    .X(\AuI.pe._092_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._534_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._085_ ),
    .B1(\AuI.pe._088_ ),
    .B2(\AuI.pe._092_ ),
    .X(\AuI.pe.Significand[7] ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._535_  (.A1(\AuI.pe._045_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._056_ ),
    .X(\AuI.pe._093_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._536_  (.A1(\AuI.pe._029_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._093_ ),
    .X(\AuI.pe._094_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._537_  (.A(\AuI.pe.significand[15] ),
    .Y(\AuI.pe._095_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._538_  (.A(\AuI.pe._095_ ),
    .B(\AuI.pe._370_ ),
    .Y(\AuI.pe._096_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._539_  (.A(\AuI.pe._096_ ),
    .X(\AuI.pe._097_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._540_  (.A1(\AuI.pe._393_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._023_ ),
    .B2(\AuI.pe.significand[7] ),
    .C1(\AuI.pe._037_ ),
    .X(\AuI.pe._098_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._541_  (.A1(\AuI.pe._062_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._072_ ),
    .C1(\AuI.pe._098_ ),
    .X(\AuI.pe._099_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._542_  (.A1(\AuI.pe._055_ ),
    .A2(\AuI.pe._079_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._020_ ),
    .C1(\AuI.pe._099_ ),
    .X(\AuI.pe._100_ ));
 sky130_fd_sc_hd__or3_4 \AuI.pe._543_  (.A(\AuI.pe.significand[8] ),
    .B(\AuI.pe._375_ ),
    .C(\AuI.pe._049_ ),
    .X(\AuI.pe._101_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._544_  (.A(\AuI.pe._393_ ),
    .X(\AuI.pe._102_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._545_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._070_ ),
    .B1(\AuI.pe._102_ ),
    .Y(\AuI.pe._103_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._546_  (.A1(\AuI.pe._101_ ),
    .A2(\AuI.pe._103_ ),
    .B1(\AuI.pe._074_ ),
    .X(\AuI.pe._104_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._547_  (.A1(\AuI.pe._094_ ),
    .A2(\AuI.pe._100_ ),
    .B1(\AuI.pe._104_ ),
    .X(\AuI.pe.Significand[8] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._548_  (.A(\AuI.pe.significand[9] ),
    .X(\AuI.pe._105_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._549_  (.A(\AuI.pe._105_ ),
    .X(\AuI.pe._106_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._550_  (.A(\AuI.pe._106_ ),
    .B(\AuI.pe._101_ ),
    .Y(\AuI.pe._107_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._551_  (.A(\AuI.pe._106_ ),
    .B(\AuI.pe._101_ ),
    .Y(\AuI.pe._108_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._552_  (.A_N(\AuI.pe._107_ ),
    .B(\AuI.pe._108_ ),
    .X(\AuI.pe._109_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._553_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._063_ ),
    .X(\AuI.pe._110_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._554_  (.A1(\AuI.pe._055_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._110_ ),
    .X(\AuI.pe._111_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._555_  (.A(\AuI.pe._391_ ),
    .X(\AuI.pe._112_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._556_  (.A1(\AuI.pe._105_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._113_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._557_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._023_ ),
    .B2(\AuI.pe._393_ ),
    .C1(\AuI.pe._113_ ),
    .X(\AuI.pe._114_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._558_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._042_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._013_ ),
    .C1(\AuI.pe._114_ ),
    .X(\AuI.pe._115_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._559_  (.A1(\AuI.pe._030_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._079_ ),
    .B2(\AuI.pe._046_ ),
    .C1(\AuI.pe._115_ ),
    .X(\AuI.pe._116_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._560_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._109_ ),
    .B1(\AuI.pe._111_ ),
    .B2(\AuI.pe._116_ ),
    .X(\AuI.pe.Significand[9] ));
 sky130_fd_sc_hd__nor3_1 \AuI.pe._561_  (.A(\AuI.pe.significand[14] ),
    .B(\AuI.pe.significand[15] ),
    .C(\AuI.pe._367_ ),
    .Y(\AuI.pe._117_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._562_  (.A(\AuI.pe.significand[13] ),
    .B(\AuI.pe._383_ ),
    .C(\AuI.pe._387_ ),
    .D(\AuI.pe._117_ ),
    .X(\AuI.pe._118_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._563_  (.A(\AuI.pe._118_ ),
    .X(\AuI.pe._119_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._564_  (.A(\AuI.pe.significand[15] ),
    .X(\AuI.pe._120_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._565_  (.A(\AuI.pe._033_ ),
    .B(\AuI.pe._120_ ),
    .C(\AuI.pe._388_ ),
    .X(\AuI.pe._121_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._566_  (.A1(\AuI.pe._028_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe._030_ ),
    .C1(\AuI.pe._121_ ),
    .X(\AuI.pe._122_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._567_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._072_ ),
    .X(\AuI.pe._123_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._568_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._123_ ),
    .X(\AuI.pe._124_ ));
 sky130_fd_sc_hd__clkbuf_4 \AuI.pe._569_  (.A(\AuI.pe._380_ ),
    .X(\AuI.pe._125_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._570_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._037_ ),
    .X(\AuI.pe._126_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._571_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._023_ ),
    .B1(\AuI.pe._042_ ),
    .B2(\AuI.pe._102_ ),
    .C1(\AuI.pe._126_ ),
    .X(\AuI.pe._127_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._572_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._079_ ),
    .B2(\AuI.pe._059_ ),
    .C1(\AuI.pe._127_ ),
    .X(\AuI.pe._128_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._573_  (.A(\AuI.pe._125_ ),
    .B(\AuI.pe._107_ ),
    .Y(\AuI.pe._129_ ));
 sky130_fd_sc_hd__o32a_1 \AuI.pe._574_  (.A1(\AuI.pe._122_ ),
    .A2(\AuI.pe._124_ ),
    .A3(\AuI.pe._128_ ),
    .B1(\AuI.pe._129_ ),
    .B2(\AuI.pe._074_ ),
    .X(\AuI.pe.Significand[10] ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._575_  (.A(\AuI.pe._028_ ),
    .B(\AuI.pe._119_ ),
    .X(\AuI.pe._130_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._576_  (.A1(\AuI.pe._055_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._046_ ),
    .C1(\AuI.pe._130_ ),
    .X(\AuI.pe._131_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._577_  (.A(\AuI.pe.significand[12] ),
    .B(\AuI.pe._388_ ),
    .C(\AuI.pe._389_ ),
    .X(\AuI.pe._132_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._578_  (.A(\AuI.pe._132_ ),
    .X(\AuI.pe._133_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._579_  (.A1(\AuI.pe._378_ ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._037_ ),
    .X(\AuI.pe._134_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._580_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._022_ ),
    .B1(\AuI.pe._041_ ),
    .B2(\AuI.pe._105_ ),
    .C1(\AuI.pe._134_ ),
    .X(\AuI.pe._135_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._581_  (.A1(\AuI.pe._102_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._079_ ),
    .B2(\AuI.pe._063_ ),
    .C1(\AuI.pe._135_ ),
    .X(\AuI.pe._136_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._582_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._089_ ),
    .X(\AuI.pe._137_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._583_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._137_ ),
    .X(\AuI.pe._138_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._584_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._136_ ),
    .C1(\AuI.pe._138_ ),
    .X(\AuI.pe._139_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._585_  (.A(\AuI.pe._373_ ),
    .B(\AuI.pe._101_ ),
    .X(\AuI.pe._140_ ));
 sky130_fd_sc_hd__clkbuf_2 \AuI.pe._586_  (.A(\AuI.pe._140_ ),
    .X(\AuI.pe._141_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._587_  (.A(\AuI.pe._378_ ),
    .X(\AuI.pe._142_ ));
 sky130_fd_sc_hd__o31ai_1 \AuI.pe._588_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._125_ ),
    .A3(\AuI.pe._101_ ),
    .B1(\AuI.pe._142_ ),
    .Y(\AuI.pe._143_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._589_  (.A1(\AuI.pe._141_ ),
    .A2(\AuI.pe._143_ ),
    .B1(\AuI.pe._074_ ),
    .X(\AuI.pe._144_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._590_  (.A1(\AuI.pe._131_ ),
    .A2(\AuI.pe._139_ ),
    .B1(\AuI.pe._144_ ),
    .X(\AuI.pe.Significand[11] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._591_  (.A(\AuI.pe.significand[12] ),
    .X(\AuI.pe._145_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._592_  (.A(\AuI.pe._145_ ),
    .B(\AuI.pe._141_ ),
    .Y(\AuI.pe._146_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._593_  (.A(\AuI.pe._072_ ),
    .B(\AuI.pe._079_ ),
    .X(\AuI.pe._147_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._594_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._059_ ),
    .C1(\AuI.pe._147_ ),
    .X(\AuI.pe._148_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._595_  (.A(\AuI.pe._378_ ),
    .Y(\AuI.pe._149_ ));
 sky130_fd_sc_hd__nor2_4 \AuI.pe._596_  (.A(\AuI.pe._149_ ),
    .B(\AuI.pe._379_ ),
    .Y(\AuI.pe._150_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._597_  (.A1(\AuI.pe._062_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._066_ ),
    .B2(\AuI.pe._089_ ),
    .X(\AuI.pe._151_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._598_  (.A1(\AuI.pe.significand[12] ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._152_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._599_  (.A1(\AuI.pe._105_ ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._022_ ),
    .B2(\AuI.pe._378_ ),
    .C1(\AuI.pe._152_ ),
    .X(\AuI.pe._153_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._600_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._041_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe.significand[2] ),
    .C1(\AuI.pe._153_ ),
    .X(\AuI.pe._154_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._601_  (.A1(\AuI.pe._102_ ),
    .A2(\AuI.pe._054_ ),
    .B1(\AuI.pe._151_ ),
    .C1(\AuI.pe._154_ ),
    .X(\AuI.pe._155_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._602_  (.A1(\AuI.pe._029_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._150_ ),
    .B2(\AuI.pe._030_ ),
    .C1(\AuI.pe._155_ ),
    .X(\AuI.pe._156_ ));
 sky130_fd_sc_hd__o2bb2a_1 \AuI.pe._603_  (.A1_N(\AuI.pe._037_ ),
    .A2_N(\AuI.pe._146_ ),
    .B1(\AuI.pe._148_ ),
    .B2(\AuI.pe._156_ ),
    .X(\AuI.pe.Significand[12] ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._604_  (.A1(\AuI.pe._102_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._054_ ),
    .B2(\AuI.pe._106_ ),
    .X(\AuI.pe._157_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._605_  (.A(\AuI.pe.significand[13] ),
    .X(\AuI.pe._158_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._606_  (.A1(\AuI.pe._158_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._159_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._607_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._022_ ),
    .B1(\AuI.pe._041_ ),
    .B2(\AuI.pe._142_ ),
    .C1(\AuI.pe._159_ ),
    .X(\AuI.pe._160_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._608_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._078_ ),
    .B2(\AuI.pe._089_ ),
    .C1(\AuI.pe._160_ ),
    .X(\AuI.pe._161_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._609_  (.A1(\AuI.pe._072_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._157_ ),
    .C1(\AuI.pe._161_ ),
    .X(\AuI.pe._162_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._610_  (.A1(\AuI.pe._055_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._150_ ),
    .B2(\AuI.pe._029_ ),
    .X(\AuI.pe._163_ ));
 sky130_fd_sc_hd__and3_2 \AuI.pe._611_  (.A(\AuI.pe._380_ ),
    .B(\AuI.pe._149_ ),
    .C(\AuI.pe._395_ ),
    .X(\AuI.pe._164_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._612_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._097_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe._045_ ),
    .X(\AuI.pe._165_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._613_  (.A1(\AuI.pe._030_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._112_ ),
    .B2(\AuI.pe._059_ ),
    .C1(\AuI.pe._165_ ),
    .X(\AuI.pe._166_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._614_  (.A(\AuI.pe._145_ ),
    .B(\AuI.pe._158_ ),
    .C(\AuI.pe._141_ ),
    .X(\AuI.pe._167_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._615_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._141_ ),
    .B1(\AuI.pe._158_ ),
    .Y(\AuI.pe._168_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._616_  (.A1(\AuI.pe._167_ ),
    .A2(\AuI.pe._168_ ),
    .B1(\AuI.pe._024_ ),
    .X(\AuI.pe._169_ ));
 sky130_fd_sc_hd__o31a_1 \AuI.pe._617_  (.A1(\AuI.pe._162_ ),
    .A2(\AuI.pe._163_ ),
    .A3(\AuI.pe._166_ ),
    .B1(\AuI.pe._169_ ),
    .X(\AuI.pe.Significand[13] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._618_  (.A(\AuI.pe.significand[14] ),
    .X(\AuI.pe._170_ ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._619_  (.A(\AuI.pe._170_ ),
    .B(\AuI.pe._167_ ),
    .X(\AuI.pe._171_ ));
 sky130_fd_sc_hd__and4b_1 \AuI.pe._620_  (.A_N(\AuI.pe.significand[10] ),
    .B(\AuI.pe._149_ ),
    .C(\AuI.pe._395_ ),
    .D(\AuI.pe._105_ ),
    .X(\AuI.pe._172_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._621_  (.A(\AuI.pe._172_ ),
    .X(\AuI.pe._173_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._622_  (.A(\AuI.pe._033_ ),
    .B(\AuI.pe._142_ ),
    .C(\AuI.pe._395_ ),
    .X(\AuI.pe._174_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._623_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._030_ ),
    .C1(\AuI.pe._174_ ),
    .X(\AuI.pe._175_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._624_  (.A(\AuI.pe.significand[4] ),
    .B(\AuI.pe._119_ ),
    .X(\AuI.pe._176_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._625_  (.A1(\AuI.pe._062_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._072_ ),
    .C1(\AuI.pe._176_ ),
    .X(\AuI.pe._177_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._626_  (.A1(\AuI.pe._089_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe._125_ ),
    .X(\AuI.pe._178_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._627_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._179_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._628_  (.A1(\AuI.pe._378_ ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._022_ ),
    .B2(\AuI.pe._158_ ),
    .C1(\AuI.pe._179_ ),
    .X(\AuI.pe._180_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._629_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._041_ ),
    .B1(\AuI.pe._078_ ),
    .B2(\AuI.pe._393_ ),
    .C1(\AuI.pe._180_ ),
    .X(\AuI.pe._181_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._630_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._066_ ),
    .B1(\AuI.pe._178_ ),
    .C1(\AuI.pe._181_ ),
    .X(\AuI.pe._182_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._631_  (.A1(\AuI.pe._029_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._177_ ),
    .C1(\AuI.pe._182_ ),
    .X(\AuI.pe._183_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._632_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._171_ ),
    .B1(\AuI.pe._175_ ),
    .B2(\AuI.pe._183_ ),
    .X(\AuI.pe.Significand[14] ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._633_  (.A(\AuI.pe._170_ ),
    .B(\AuI.pe._167_ ),
    .X(\AuI.pe._184_ ));
 sky130_fd_sc_hd__o2bb2a_1 \AuI.pe._634_  (.A1_N(\AuI.pe._120_ ),
    .A2_N(\AuI.pe._184_ ),
    .B1(\AuI.pe._141_ ),
    .B2(\AuI.pe._372_ ),
    .X(\AuI.pe._185_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._635_  (.A(\AuI.pe._045_ ),
    .B(\AuI.pe._142_ ),
    .C(\AuI.pe._395_ ),
    .X(\AuI.pe._186_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._636_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._029_ ),
    .C1(\AuI.pe._186_ ),
    .X(\AuI.pe._187_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._637_  (.A1(\AuI.pe._105_ ),
    .A2(\AuI.pe._078_ ),
    .B1(\AuI.pe._097_ ),
    .B2(\AuI.pe._089_ ),
    .X(\AuI.pe._188_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._638_  (.A1(\AuI.pe._393_ ),
    .A2(\AuI.pe._399_ ),
    .B1(\AuI.pe._002_ ),
    .B2(\AuI.pe._380_ ),
    .X(\AuI.pe._189_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._639_  (.A1(\AuI.pe._120_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._190_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._640_  (.A1(\AuI.pe.significand[12] ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._022_ ),
    .B2(\AuI.pe._170_ ),
    .C1(\AuI.pe._190_ ),
    .X(\AuI.pe._191_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._641_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._391_ ),
    .B1(\AuI.pe._041_ ),
    .B2(\AuI.pe._158_ ),
    .C1(\AuI.pe._191_ ),
    .X(\AuI.pe._192_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._642_  (.A1(\AuI.pe._142_ ),
    .A2(\AuI.pe._053_ ),
    .B1(\AuI.pe._189_ ),
    .C1(\AuI.pe._192_ ),
    .X(\AuI.pe._193_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._643_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._119_ ),
    .B1(\AuI.pe._188_ ),
    .C1(\AuI.pe._193_ ),
    .X(\AuI.pe._194_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._644_  (.A1(\AuI.pe._055_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._397_ ),
    .B2(\AuI.pe._030_ ),
    .C1(\AuI.pe._194_ ),
    .X(\AuI.pe._195_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._645_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._185_ ),
    .B1(\AuI.pe._187_ ),
    .B2(\AuI.pe._195_ ),
    .X(\AuI.pe.Significand[15] ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._646_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._055_ ),
    .X(\AuI.pe._196_ ));
 sky130_fd_sc_hd__nor2_4 \AuI.pe._647_  (.A(\AuI.pe._370_ ),
    .B(\AuI.pe._374_ ),
    .Y(\AuI.pe._197_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._648_  (.A1(\AuI.pe._030_ ),
    .A2(\AuI.pe._084_ ),
    .A3(\AuI.pe._197_ ),
    .B1(\AuI.pe._150_ ),
    .B2(\AuI.pe._059_ ),
    .X(\AuI.pe._198_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._649_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._078_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe._071_ ),
    .X(\AuI.pe._199_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._650_  (.A1(\AuI.pe._378_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe.significand[12] ),
    .X(\AuI.pe._200_ ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._651_  (.A(\AuI.pe._367_ ),
    .X(\AuI.pe._201_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._652_  (.A1(\AuI.pe._201_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._036_ ),
    .X(\AuI.pe._202_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._653_  (.A1(\AuI.pe.significand[13] ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._006_ ),
    .B2(\AuI.pe._120_ ),
    .C1(\AuI.pe._202_ ),
    .X(\AuI.pe._203_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._654_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._041_ ),
    .B1(\AuI.pe._096_ ),
    .B2(\AuI.pe._393_ ),
    .C1(\AuI.pe._203_ ),
    .X(\AuI.pe._204_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._655_  (.A1(\AuI.pe._105_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._200_ ),
    .C1(\AuI.pe._204_ ),
    .X(\AuI.pe._205_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._656_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._199_ ),
    .C1(\AuI.pe._205_ ),
    .X(\AuI.pe._206_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._657_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._397_ ),
    .B2(\AuI.pe._028_ ),
    .C1(\AuI.pe._206_ ),
    .X(\AuI.pe._207_ ));
 sky130_fd_sc_hd__or4_2 \AuI.pe._658_  (.A(\AuI.pe._201_ ),
    .B(\AuI.pe._372_ ),
    .C(\AuI.pe._373_ ),
    .D(\AuI.pe._101_ ),
    .X(\AuI.pe._208_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._659_  (.A1(\AuI.pe._372_ ),
    .A2(\AuI.pe._141_ ),
    .B1(\AuI.pe._201_ ),
    .Y(\AuI.pe._209_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._660_  (.A1(\AuI.pe._208_ ),
    .A2(\AuI.pe._209_ ),
    .B1(\AuI.pe._024_ ),
    .X(\AuI.pe._210_ ));
 sky130_fd_sc_hd__o31a_1 \AuI.pe._661_  (.A1(\AuI.pe._196_ ),
    .A2(\AuI.pe._198_ ),
    .A3(\AuI.pe._207_ ),
    .B1(\AuI.pe._210_ ),
    .X(\AuI.pe.Significand[16] ));
 sky130_fd_sc_hd__buf_2 \AuI.pe._662_  (.A(\AuI.pe.significand[17] ),
    .X(\AuI.pe._211_ ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._663_  (.A(\AuI.pe._211_ ),
    .B(\AuI.pe._208_ ),
    .X(\AuI.pe._212_ ));
 sky130_fd_sc_hd__and3b_2 \AuI.pe._664_  (.A_N(\AuI.pe.significand[7] ),
    .B(\AuI.pe._197_ ),
    .C(\AuI.pe._071_ ),
    .X(\AuI.pe._213_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._665_  (.A1(\AuI.pe._033_ ),
    .A2(\AuI.pe._397_ ),
    .B1(\AuI.pe._213_ ),
    .B2(\AuI.pe._014_ ),
    .X(\AuI.pe._214_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._666_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._214_ ),
    .X(\AuI.pe._215_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._667_  (.A1(\AuI.pe._013_ ),
    .A2(\AuI.pe.significand[7] ),
    .A3(\AuI.pe._197_ ),
    .B1(\AuI.pe._150_ ),
    .B2(\AuI.pe._062_ ),
    .X(\AuI.pe._216_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._668_  (.A1(\AuI.pe._072_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._045_ ),
    .C1(\AuI.pe._216_ ),
    .X(\AuI.pe._217_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._669_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._384_ ),
    .A3(\AuI.pe._387_ ),
    .B1(\AuI.pe._023_ ),
    .X(\AuI.pe._218_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._670_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._119_ ),
    .B1(\AuI.pe._218_ ),
    .B2(\AuI.pe._201_ ),
    .X(\AuI.pe._219_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._671_  (.A1(\AuI.pe._211_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._041_ ),
    .B2(\AuI.pe._120_ ),
    .C1(\AuI.pe._036_ ),
    .X(\AuI.pe._220_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._672_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe._158_ ),
    .X(\AuI.pe._221_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._673_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._050_ ),
    .B1(\AuI.pe._220_ ),
    .C1(\AuI.pe._221_ ),
    .X(\AuI.pe._222_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._674_  (.A1(\AuI.pe._102_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._079_ ),
    .B2(\AuI.pe._142_ ),
    .C1(\AuI.pe._222_ ),
    .X(\AuI.pe._223_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI.pe._675_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._097_ ),
    .B1(\AuI.pe._217_ ),
    .C1(\AuI.pe._219_ ),
    .D1(\AuI.pe._223_ ),
    .X(\AuI.pe._224_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._676_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._212_ ),
    .B1(\AuI.pe._215_ ),
    .B2(\AuI.pe._224_ ),
    .X(\AuI.pe.Significand[17] ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._677_  (.A(\AuI.pe._062_ ),
    .B(\AuI.pe._197_ ),
    .C(\AuI.pe._010_ ),
    .X(\AuI.pe._225_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._678_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._213_ ),
    .B2(\AuI.pe._028_ ),
    .X(\AuI.pe._226_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._679_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._397_ ),
    .B1(\AuI.pe._225_ ),
    .B2(\AuI.pe._030_ ),
    .C1(\AuI.pe._226_ ),
    .X(\AuI.pe._227_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._680_  (.A(\AuI.pe.significand[2] ),
    .B(\AuI.pe.significand[7] ),
    .C(\AuI.pe._197_ ),
    .X(\AuI.pe._228_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._681_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._150_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe.significand[4] ),
    .X(\AuI.pe._229_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._682_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._228_ ),
    .C1(\AuI.pe._229_ ),
    .X(\AuI.pe._230_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._683_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._079_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe._102_ ),
    .X(\AuI.pe._231_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._684_  (.A1(\AuI.pe._158_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe._170_ ),
    .X(\AuI.pe._232_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._685_  (.A1(\AuI.pe._142_ ),
    .A2(\AuI.pe._086_ ),
    .B1(\AuI.pe._232_ ),
    .X(\AuI.pe._233_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._686_  (.A1(\AuI.pe._385_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._022_ ),
    .B2(\AuI.pe._211_ ),
    .C1(\AuI.pe._036_ ),
    .X(\AuI.pe._234_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._687_  (.A1(\AuI.pe._120_ ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._041_ ),
    .B2(\AuI.pe._201_ ),
    .C1(\AuI.pe._234_ ),
    .X(\AuI.pe._235_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._688_  (.A1(\AuI.pe._125_ ),
    .A2(\AuI.pe._097_ ),
    .B1(\AuI.pe._233_ ),
    .C1(\AuI.pe._235_ ),
    .X(\AuI.pe._236_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI.pe._689_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._230_ ),
    .C1(\AuI.pe._231_ ),
    .D1(\AuI.pe._236_ ),
    .X(\AuI.pe._237_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._690_  (.A(\AuI.pe._211_ ),
    .B(\AuI.pe._385_ ),
    .C(\AuI.pe._208_ ),
    .X(\AuI.pe._238_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._691_  (.A1(\AuI.pe._211_ ),
    .A2(\AuI.pe._208_ ),
    .B1(\AuI.pe._385_ ),
    .Y(\AuI.pe._239_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._692_  (.A1(\AuI.pe._238_ ),
    .A2(\AuI.pe._239_ ),
    .B1(\AuI.pe._024_ ),
    .X(\AuI.pe._240_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._693_  (.A1(\AuI.pe._227_ ),
    .A2(\AuI.pe._237_ ),
    .B1(\AuI.pe._240_ ),
    .X(\AuI.pe.Significand[18] ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._694_  (.A(\AuI.pe._386_ ),
    .B(\AuI.pe._238_ ),
    .X(\AuI.pe._241_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._695_  (.A(\AuI.pe._014_ ),
    .B(\AuI.pe._012_ ),
    .X(\AuI.pe._242_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._696_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._397_ ),
    .B1(\AuI.pe._213_ ),
    .B2(\AuI.pe._055_ ),
    .C1(\AuI.pe._242_ ),
    .X(\AuI.pe._243_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._697_  (.A1(\AuI.pe._089_ ),
    .A2(\AuI.pe._150_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._062_ ),
    .X(\AuI.pe._244_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._698_  (.A1(\AuI.pe._045_ ),
    .A2(\AuI.pe._089_ ),
    .A3(\AuI.pe._197_ ),
    .B1(\AuI.pe._133_ ),
    .B2(\AuI.pe._102_ ),
    .X(\AuI.pe._245_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._699_  (.A1(\AuI.pe._380_ ),
    .A2(\AuI.pe._391_ ),
    .B1(\AuI.pe._118_ ),
    .B2(\AuI.pe._105_ ),
    .X(\AuI.pe._246_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._700_  (.A1(\AuI.pe._386_ ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe._078_ ),
    .B2(\AuI.pe.significand[13] ),
    .C1(\AuI.pe._036_ ),
    .X(\AuI.pe._247_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._701_  (.A1(\AuI.pe._201_ ),
    .A2(\AuI.pe._004_ ),
    .B1(\AuI.pe._040_ ),
    .B2(\AuI.pe._211_ ),
    .X(\AuI.pe._248_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._702_  (.A1(\AuI.pe._385_ ),
    .A2(\AuI.pe._022_ ),
    .B1(\AuI.pe._247_ ),
    .C1(\AuI.pe._248_ ),
    .X(\AuI.pe._249_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._703_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe._120_ ),
    .X(\AuI.pe._250_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._704_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._399_ ),
    .B1(\AuI.pe._249_ ),
    .C1(\AuI.pe._250_ ),
    .X(\AuI.pe._251_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._705_  (.A1(\AuI.pe._142_ ),
    .A2(\AuI.pe._097_ ),
    .B1(\AuI.pe._246_ ),
    .C1(\AuI.pe._251_ ),
    .X(\AuI.pe._252_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._706_  (.A1(\AuI.pe._072_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._225_ ),
    .B2(\AuI.pe._013_ ),
    .X(\AuI.pe._253_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._707_  (.A(\AuI.pe._244_ ),
    .B(\AuI.pe._245_ ),
    .C(\AuI.pe._252_ ),
    .D(\AuI.pe._253_ ),
    .X(\AuI.pe._254_ ));
 sky130_fd_sc_hd__o22a_1 \AuI.pe._708_  (.A1(\AuI.pe._074_ ),
    .A2(\AuI.pe._241_ ),
    .B1(\AuI.pe._243_ ),
    .B2(\AuI.pe._254_ ),
    .X(\AuI.pe.Significand[19] ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._709_  (.A(\AuI.pe._393_ ),
    .B(\AuI.pe._375_ ),
    .Y(\AuI.pe._255_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._710_  (.A(\AuI.pe.significand[3] ),
    .B(\AuI.pe._394_ ),
    .C(\AuI.pe._395_ ),
    .D(\AuI.pe._255_ ),
    .X(\AuI.pe._256_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._711_  (.A1(\AuI.pe._063_ ),
    .A2(\AuI.pe._397_ ),
    .B1(\AuI.pe._256_ ),
    .B2(\AuI.pe._014_ ),
    .X(\AuI.pe._257_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._712_  (.A1(\AuI.pe._084_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._225_ ),
    .B2(\AuI.pe._055_ ),
    .C1(\AuI.pe._257_ ),
    .X(\AuI.pe._258_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._713_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._089_ ),
    .A3(\AuI.pe._197_ ),
    .B1(\AuI.pe._150_ ),
    .B2(\AuI.pe._102_ ),
    .X(\AuI.pe._259_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._714_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._133_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._071_ ),
    .X(\AuI.pe._260_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._715_  (.A1(\AuI.pe._145_ ),
    .A2(\AuI.pe._096_ ),
    .B1(\AuI.pe._118_ ),
    .B2(\AuI.pe._380_ ),
    .X(\AuI.pe._261_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._716_  (.A1(\AuI.pe.significand[20] ),
    .A2(\AuI.pe.significand[23] ),
    .B1(\AuI.pe._035_ ),
    .X(\AuI.pe._262_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._717_  (.A1(\AuI.pe._386_ ),
    .A2(\AuI.pe._006_ ),
    .B1(\AuI.pe._040_ ),
    .B2(\AuI.pe._385_ ),
    .C1(\AuI.pe._262_ ),
    .X(\AuI.pe._263_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._718_  (.A1(\AuI.pe._120_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._004_ ),
    .B2(\AuI.pe._211_ ),
    .C1(\AuI.pe._263_ ),
    .X(\AuI.pe._264_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._719_  (.A1(\AuI.pe._158_ ),
    .A2(\AuI.pe._399_ ),
    .B1(\AuI.pe._053_ ),
    .B2(\AuI.pe._201_ ),
    .X(\AuI.pe._265_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._720_  (.A1(\AuI.pe._142_ ),
    .A2(\AuI.pe._112_ ),
    .B1(\AuI.pe._264_ ),
    .C1(\AuI.pe._265_ ),
    .X(\AuI.pe._266_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._721_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._078_ ),
    .B1(\AuI.pe._261_ ),
    .C1(\AuI.pe._266_ ),
    .X(\AuI.pe._267_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._722_  (.A1(\AuI.pe._013_ ),
    .A2(\AuI.pe._012_ ),
    .B1(\AuI.pe._213_ ),
    .B2(\AuI.pe._045_ ),
    .X(\AuI.pe._268_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._723_  (.A(\AuI.pe._259_ ),
    .B(\AuI.pe._260_ ),
    .C(\AuI.pe._267_ ),
    .D(\AuI.pe._268_ ),
    .X(\AuI.pe._269_ ));
 sky130_fd_sc_hd__or4b_1 \AuI.pe._724_  (.A(\AuI.pe._211_ ),
    .B(\AuI.pe._208_ ),
    .C(\AuI.pe.significand[20] ),
    .D_N(\AuI.pe._076_ ),
    .X(\AuI.pe._270_ ));
 sky130_fd_sc_hd__o21ai_1 \AuI.pe._725_  (.A1(\AuI.pe._386_ ),
    .A2(\AuI.pe._238_ ),
    .B1(\AuI.pe.significand[20] ),
    .Y(\AuI.pe._271_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._726_  (.A1(\AuI.pe._270_ ),
    .A2(\AuI.pe._271_ ),
    .B1(\AuI.pe._024_ ),
    .X(\AuI.pe._272_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._727_  (.A1(\AuI.pe._258_ ),
    .A2(\AuI.pe._269_ ),
    .B1(\AuI.pe._272_ ),
    .X(\AuI.pe.Significand[20] ));
 sky130_fd_sc_hd__nand2_2 \AuI.pe._728_  (.A(\AuI.pe._388_ ),
    .B(\AuI.pe._009_ ),
    .Y(\AuI.pe._273_ ));
 sky130_fd_sc_hd__nor3_1 \AuI.pe._729_  (.A(\AuI.pe._273_ ),
    .B(\AuI.pe._375_ ),
    .C(\AuI.pe._376_ ),
    .Y(\AuI.pe._274_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._730_  (.A1(\AuI.pe._033_ ),
    .A2(\AuI.pe._012_ ),
    .B1(\AuI.pe._256_ ),
    .B2(\AuI.pe._028_ ),
    .X(\AuI.pe._275_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._731_  (.A1(\AuI.pe._020_ ),
    .A2(\AuI.pe._274_ ),
    .B1(\AuI.pe._275_ ),
    .X(\AuI.pe._276_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._732_  (.A1(\AuI.pe._062_ ),
    .A2(\AuI.pe._197_ ),
    .B1(\AuI.pe._173_ ),
    .X(\AuI.pe._277_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._733_  (.A1(\AuI.pe._102_ ),
    .A2(\AuI.pe._164_ ),
    .B1(\AuI.pe._397_ ),
    .B2(\AuI.pe._072_ ),
    .X(\AuI.pe._278_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._734_  (.A1(\AuI.pe._046_ ),
    .A2(\AuI.pe._225_ ),
    .B1(\AuI.pe._277_ ),
    .B2(\AuI.pe._084_ ),
    .C1(\AuI.pe._278_ ),
    .X(\AuI.pe._279_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._735_  (.A1(\AuI.pe.significand[21] ),
    .A2(\AuI.pe._026_ ),
    .B1(\AuI.pe._002_ ),
    .B2(\AuI.pe._201_ ),
    .C1(\AuI.pe._037_ ),
    .X(\AuI.pe._280_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._736_  (.A1(\AuI.pe._385_ ),
    .A2(\AuI.pe._384_ ),
    .B1(\AuI.pe._022_ ),
    .X(\AuI.pe._281_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._737_  (.A1(\AuI.pe._170_ ),
    .A2(\AuI.pe._399_ ),
    .B1(\AuI.pe._281_ ),
    .B2(\AuI.pe.significand[20] ),
    .X(\AuI.pe._282_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._738_  (.A1(\AuI.pe._158_ ),
    .A2(\AuI.pe._096_ ),
    .B1(\AuI.pe._119_ ),
    .B2(\AuI.pe._142_ ),
    .X(\AuI.pe._283_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI.pe._739_  (.A1(\AuI.pe._106_ ),
    .A2(\AuI.pe._150_ ),
    .B1(\AuI.pe._280_ ),
    .C1(\AuI.pe._282_ ),
    .D1(\AuI.pe._283_ ),
    .X(\AuI.pe._284_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._740_  (.A1(\AuI.pe._211_ ),
    .A2(\AuI.pe._000_ ),
    .A3(\AuI.pe._384_ ),
    .B1(\AuI.pe._042_ ),
    .X(\AuI.pe._285_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._741_  (.A1(\AuI.pe._380_ ),
    .A2(\AuI.pe._389_ ),
    .B1(\AuI.pe._390_ ),
    .X(\AuI.pe._286_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._742_  (.A(\AuI.pe._145_ ),
    .B(\AuI.pe._388_ ),
    .C(\AuI.pe._286_ ),
    .X(\AuI.pe._287_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._743_  (.A1(\AuI.pe._120_ ),
    .A2(\AuI.pe._079_ ),
    .B1(\AuI.pe._285_ ),
    .B2(\AuI.pe._386_ ),
    .C1(\AuI.pe._287_ ),
    .X(\AuI.pe._288_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._744_  (.A1(\AuI.pe._059_ ),
    .A2(\AuI.pe._213_ ),
    .B1(\AuI.pe._284_ ),
    .C1(\AuI.pe._288_ ),
    .X(\AuI.pe._289_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._745_  (.A(\AuI.pe.significand[21] ),
    .B(\AuI.pe._270_ ),
    .Y(\AuI.pe._290_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._746_  (.A(\AuI.pe.significand[21] ),
    .B(\AuI.pe._270_ ),
    .X(\AuI.pe._291_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._747_  (.A1(\AuI.pe._290_ ),
    .A2(\AuI.pe._291_ ),
    .B1(\AuI.pe._024_ ),
    .X(\AuI.pe._292_ ));
 sky130_fd_sc_hd__o31a_1 \AuI.pe._748_  (.A1(\AuI.pe._276_ ),
    .A2(\AuI.pe._279_ ),
    .A3(\AuI.pe._289_ ),
    .B1(\AuI.pe._292_ ),
    .X(\AuI.pe.Significand[21] ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._749_  (.A(\AuI.pe.significand[22] ),
    .B(\AuI.pe._291_ ),
    .Y(\AuI.pe._293_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._750_  (.A(\AuI.pe._024_ ),
    .B(\AuI.pe._293_ ),
    .X(\AuI.pe._294_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._751_  (.A1(\AuI.pe.significand[22] ),
    .A2(\AuI.pe._291_ ),
    .B1(\AuI.pe._294_ ),
    .Y(\AuI.pe._295_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._752_  (.A1(\AuI.pe._013_ ),
    .A2(\AuI.pe._274_ ),
    .B1(\AuI.pe._256_ ),
    .B2(\AuI.pe.significand[2] ),
    .X(\AuI.pe._296_ ));
 sky130_fd_sc_hd__or3b_1 \AuI.pe._753_  (.A(\AuI.pe.significand[2] ),
    .B(\AuI.pe.significand[3] ),
    .C_N(\AuI.pe._013_ ),
    .X(\AuI.pe._297_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._754_  (.A(\AuI.pe.significand[8] ),
    .B(\AuI.pe._375_ ),
    .C(\AuI.pe._297_ ),
    .X(\AuI.pe._298_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._755_  (.A(\AuI.pe._373_ ),
    .B(\AuI.pe._379_ ),
    .C(\AuI.pe._298_ ),
    .X(\AuI.pe._299_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._756_  (.A(\AuI.pe._299_ ),
    .Y(\AuI.pe._300_ ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._757_  (.A1(\AuI.pe._158_ ),
    .A2(\AuI.pe._391_ ),
    .B1(\AuI.pe._118_ ),
    .B2(\AuI.pe.significand[12] ),
    .X(\AuI.pe._301_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._758_  (.A1(\AuI.pe.significand[5] ),
    .A2(\AuI.pe._213_ ),
    .B1(\AuI.pe._078_ ),
    .B2(\AuI.pe._201_ ),
    .C1(\AuI.pe._301_ ),
    .X(\AuI.pe._302_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._759_  (.A1(\AuI.pe.significand[3] ),
    .A2(\AuI.pe._012_ ),
    .B1(\AuI.pe._300_ ),
    .B2(\AuI.pe._014_ ),
    .C1(\AuI.pe._302_ ),
    .X(\AuI.pe._303_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._760_  (.A1(\AuI.pe._071_ ),
    .A2(\AuI.pe._197_ ),
    .B1(\AuI.pe._397_ ),
    .X(\AuI.pe._304_ ));
 sky130_fd_sc_hd__o211a_1 \AuI.pe._761_  (.A1(\AuI.pe._385_ ),
    .A2(\AuI.pe.significand[20] ),
    .B1(\AuI.pe._384_ ),
    .C1(\AuI.pe._386_ ),
    .X(\AuI.pe._305_ ));
 sky130_fd_sc_hd__o211a_1 \AuI.pe._762_  (.A1(\AuI.pe.significand[21] ),
    .A2(\AuI.pe._025_ ),
    .B1(\AuI.pe.significand[22] ),
    .C1(\AuI.pe.significand[24] ),
    .X(\AuI.pe._306_ ));
 sky130_fd_sc_hd__o2111a_1 \AuI.pe._763_  (.A1(\AuI.pe.significand[14] ),
    .A2(\AuI.pe._201_ ),
    .B1(\AuI.pe._384_ ),
    .C1(\AuI.pe._387_ ),
    .D1(\AuI.pe._120_ ),
    .X(\AuI.pe._307_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI.pe._764_  (.A1(\AuI.pe.significand[20] ),
    .A2(\AuI.pe._041_ ),
    .B1(\AuI.pe._305_ ),
    .C1(\AuI.pe._306_ ),
    .D1(\AuI.pe._307_ ),
    .X(\AuI.pe._308_ ));
 sky130_fd_sc_hd__a221o_1 \AuI.pe._765_  (.A1(\AuI.pe._211_ ),
    .A2(\AuI.pe._002_ ),
    .B1(\AuI.pe._173_ ),
    .B2(\AuI.pe._393_ ),
    .C1(\AuI.pe._308_ ),
    .X(\AuI.pe._309_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._766_  (.A(\AuI.pe._105_ ),
    .B(\AuI.pe._378_ ),
    .X(\AuI.pe._310_ ));
 sky130_fd_sc_hd__a32o_1 \AuI.pe._767_  (.A1(\AuI.pe._380_ ),
    .A2(\AuI.pe._395_ ),
    .A3(\AuI.pe._310_ ),
    .B1(\AuI.pe._132_ ),
    .B2(\AuI.pe._378_ ),
    .X(\AuI.pe._311_ ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._768_  (.A1(\AuI.pe._089_ ),
    .A2(\AuI.pe._304_ ),
    .B1(\AuI.pe._309_ ),
    .C1(\AuI.pe._311_ ),
    .X(\AuI.pe._312_ ));
 sky130_fd_sc_hd__a2111o_1 \AuI.pe._769_  (.A1(\AuI.pe._056_ ),
    .A2(\AuI.pe._225_ ),
    .B1(\AuI.pe._296_ ),
    .C1(\AuI.pe._303_ ),
    .D1(\AuI.pe._312_ ),
    .X(\AuI.pe._313_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._770_  (.A(\AuI.pe._295_ ),
    .B(\AuI.pe._313_ ),
    .X(\AuI.pe._314_ ));
 sky130_fd_sc_hd__clkbuf_1 \AuI.pe._771_  (.A(\AuI.pe._314_ ),
    .X(\AuI.pe.Significand[22] ));
 sky130_fd_sc_hd__a41o_1 \AuI.pe._777_  (.A1(\AuI.pe._377_ ),
    .A2(\AuI.pe._381_ ),
    .A3(\AuI.pe._398_ ),
    .A4(\AuI.pe._018_ ),
    .B1(\AuI.exp_a ),
    .X(\AuI.pe._318_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._778_  (.A(\AuI.operand_a[24] ),
    .Y(\AuI.pe._319_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._779_  (.A(\AuI.pe._399_ ),
    .B(\AuI.pe._078_ ),
    .X(\AuI.pe._320_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._780_  (.A(\AuI.pe._003_ ),
    .B(\AuI.pe._040_ ),
    .C(\AuI.pe._118_ ),
    .X(\AuI.pe._321_ ));
 sky130_fd_sc_hd__o2111a_1 \AuI.pe._781_  (.A1(\AuI.pe.significand[5] ),
    .A2(\AuI.pe.significand[4] ),
    .B1(\AuI.pe._388_ ),
    .C1(\AuI.pe._009_ ),
    .D1(\AuI.pe._010_ ),
    .X(\AuI.pe._322_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._782_  (.A(\AuI.pe._132_ ),
    .B(\AuI.pe._320_ ),
    .C(\AuI.pe._321_ ),
    .D(\AuI.pe._322_ ),
    .X(\AuI.pe._323_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._783_  (.A(\AuI.pe._016_ ),
    .B(\AuI.pe._299_ ),
    .Y(\AuI.pe._324_ ));
 sky130_fd_sc_hd__or2_1 \AuI.pe._784_  (.A(\AuI.pe._397_ ),
    .B(\AuI.pe._173_ ),
    .X(\AuI.pe._325_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._785_  (.A(\AuI.pe._319_ ),
    .B(\AuI.pe._323_ ),
    .C(\AuI.pe._324_ ),
    .D(\AuI.pe._325_ ),
    .X(\AuI.pe._326_ ));
 sky130_fd_sc_hd__o31ai_1 \AuI.pe._786_  (.A1(\AuI.pe._323_ ),
    .A2(\AuI.pe._324_ ),
    .A3(\AuI.pe._325_ ),
    .B1(\AuI.pe._319_ ),
    .Y(\AuI.pe._327_ ));
 sky130_fd_sc_hd__and3_1 \AuI.pe._787_  (.A(\AuI.pe._318_ ),
    .B(\AuI.pe._326_ ),
    .C(\AuI.pe._327_ ),
    .X(\AuI.pe._328_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._788_  (.A1(\AuI.pe._326_ ),
    .A2(\AuI.pe._327_ ),
    .B1(\AuI.pe._318_ ),
    .Y(\AuI.pe._329_ ));
 sky130_fd_sc_hd__nor2_1 \AuI.pe._789_  (.A(\AuI.pe._328_ ),
    .B(\AuI.pe._329_ ),
    .Y(\AuI.exponent_sub[1] ));
 sky130_fd_sc_hd__a21bo_1 \AuI.pe._790_  (.A1(\AuI.pe._318_ ),
    .A2(\AuI.pe._327_ ),
    .B1_N(\AuI.pe._326_ ),
    .X(\AuI.pe._330_ ));
 sky130_fd_sc_hd__and2_1 \AuI.pe._791_  (.A(\AuI.pe._016_ ),
    .B(\AuI.pe._299_ ),
    .X(\AuI.pe._331_ ));
 sky130_fd_sc_hd__o311a_1 \AuI.pe._792_  (.A1(\AuI.pe._393_ ),
    .A2(\AuI.pe._105_ ),
    .A3(\AuI.pe._380_ ),
    .B1(\AuI.pe._149_ ),
    .C1(\AuI.pe._395_ ),
    .X(\AuI.pe._332_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._793_  (.A(\AuI.pe._332_ ),
    .Y(\AuI.pe._333_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._794_  (.A(\AuI.pe.significand[20] ),
    .B(\AuI.pe._368_ ),
    .C(\AuI.pe._076_ ),
    .X(\AuI.pe._334_ ));
 sky130_fd_sc_hd__or3b_1 \AuI.pe._795_  (.A(\AuI.pe._399_ ),
    .B(\AuI.pe._078_ ),
    .C_N(\AuI.pe._334_ ),
    .X(\AuI.pe._335_ ));
 sky130_fd_sc_hd__nand2_1 \AuI.pe._796_  (.A(\AuI.pe._384_ ),
    .B(\AuI.pe._387_ ),
    .Y(\AuI.pe._336_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._797_  (.A(\AuI.pe._149_ ),
    .B(\AuI.pe._367_ ),
    .C(\AuI.pe._336_ ),
    .D(\AuI.pe._372_ ),
    .X(\AuI.pe._337_ ));
 sky130_fd_sc_hd__and4bb_1 \AuI.pe._798_  (.A_N(\AuI.pe._335_ ),
    .B_N(\AuI.pe._256_ ),
    .C(\AuI.pe._337_ ),
    .D(\AuI.pe._377_ ),
    .X(\AuI.pe._338_ ));
 sky130_fd_sc_hd__and4_1 \AuI.pe._799_  (.A(\AuI.operand_a[25] ),
    .B(\AuI.pe._331_ ),
    .C(\AuI.pe._333_ ),
    .D(\AuI.pe._338_ ),
    .X(\AuI.pe._339_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._800_  (.A1(\AuI.pe._331_ ),
    .A2(\AuI.pe._333_ ),
    .A3(\AuI.pe._338_ ),
    .B1(\AuI.operand_a[25] ),
    .X(\AuI.pe._340_ ));
 sky130_fd_sc_hd__nor2b_1 \AuI.pe._801_  (.A(\AuI.pe._339_ ),
    .B_N(\AuI.pe._340_ ),
    .Y(\AuI.pe._341_ ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._802_  (.A(\AuI.pe._330_ ),
    .B(\AuI.pe._341_ ),
    .X(\AuI.exponent_sub[2] ));
 sky130_fd_sc_hd__nor3_1 \AuI.pe._803_  (.A(\AuI.pe._273_ ),
    .B(\AuI.pe._375_ ),
    .C(\AuI.pe._049_ ),
    .Y(\AuI.pe._342_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._804_  (.A(\AuI.pe._392_ ),
    .B(\AuI.pe._096_ ),
    .C(\AuI.pe._118_ ),
    .D(\AuI.pe._150_ ),
    .X(\AuI.pe._343_ ));
 sky130_fd_sc_hd__and4bb_1 \AuI.pe._805_  (.A_N(\AuI.pe._342_ ),
    .B_N(\AuI.pe._343_ ),
    .C(\AuI.operand_a[26] ),
    .D(\AuI.pe._333_ ),
    .X(\AuI.pe._344_ ));
 sky130_fd_sc_hd__inv_2 \AuI.pe._806_  (.A(\AuI.pe._391_ ),
    .Y(\AuI.pe._345_ ));
 sky130_fd_sc_hd__clkinv_2 \AuI.pe._807_  (.A(\AuI.pe.significand[12] ),
    .Y(\AuI.pe._346_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._808_  (.A(\AuI.pe.significand[13] ),
    .B(\AuI.pe.significand[14] ),
    .C(\AuI.pe.significand[15] ),
    .D(\AuI.pe._367_ ),
    .X(\AuI.pe._347_ ));
 sky130_fd_sc_hd__or3_1 \AuI.pe._809_  (.A(\AuI.pe._346_ ),
    .B(\AuI.pe._336_ ),
    .C(\AuI.pe._347_ ),
    .X(\AuI.pe._348_ ));
 sky130_fd_sc_hd__or4b_1 \AuI.pe._810_  (.A(\AuI.pe.significand[14] ),
    .B(\AuI.pe.significand[15] ),
    .C(\AuI.pe._367_ ),
    .D_N(\AuI.pe.significand[13] ),
    .X(\AuI.pe._349_ ));
 sky130_fd_sc_hd__o221a_1 \AuI.pe._811_  (.A1(\AuI.pe._095_ ),
    .A2(\AuI.pe._370_ ),
    .B1(\AuI.pe._349_ ),
    .B2(\AuI.pe._336_ ),
    .C1(\AuI.pe._337_ ),
    .X(\AuI.pe._350_ ));
 sky130_fd_sc_hd__or4b_1 \AuI.pe._812_  (.A(\AuI.pe.significand[10] ),
    .B(\AuI.pe.significand[11] ),
    .C(\AuI.pe.significand[12] ),
    .D_N(\AuI.pe.significand[9] ),
    .X(\AuI.pe._351_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._813_  (.A(\AuI.pe._368_ ),
    .B(\AuI.pe._369_ ),
    .C(\AuI.pe._347_ ),
    .D(\AuI.pe._351_ ),
    .X(\AuI.pe._352_ ));
 sky130_fd_sc_hd__o41a_1 \AuI.pe._814_  (.A1(\AuI.pe._008_ ),
    .A2(\AuI.pe._370_ ),
    .A3(\AuI.pe._372_ ),
    .A4(\AuI.pe._373_ ),
    .B1(\AuI.pe._352_ ),
    .X(\AuI.pe._353_ ));
 sky130_fd_sc_hd__or4_1 \AuI.pe._815_  (.A(\AuI.pe._367_ ),
    .B(\AuI.pe._368_ ),
    .C(\AuI.pe._369_ ),
    .D(\AuI.pe._372_ ),
    .X(\AuI.pe._354_ ));
 sky130_fd_sc_hd__or3b_1 \AuI.pe._816_  (.A(\AuI.pe._378_ ),
    .B(\AuI.pe._354_ ),
    .C_N(\AuI.pe._380_ ),
    .X(\AuI.pe._355_ ));
 sky130_fd_sc_hd__o311a_1 \AuI.pe._817_  (.A1(\AuI.pe.significand[7] ),
    .A2(\AuI.pe._273_ ),
    .A3(\AuI.pe._070_ ),
    .B1(\AuI.pe._353_ ),
    .C1(\AuI.pe._355_ ),
    .X(\AuI.pe._356_ ));
 sky130_fd_sc_hd__a41o_1 \AuI.pe._818_  (.A1(\AuI.pe._345_ ),
    .A2(\AuI.pe._348_ ),
    .A3(\AuI.pe._350_ ),
    .A4(\AuI.pe._356_ ),
    .B1(\AuI.operand_a[26] ),
    .X(\AuI.pe._357_ ));
 sky130_fd_sc_hd__and2b_1 \AuI.pe._819_  (.A_N(\AuI.pe._344_ ),
    .B(\AuI.pe._357_ ),
    .X(\AuI.pe._358_ ));
 sky130_fd_sc_hd__a21oi_1 \AuI.pe._820_  (.A1(\AuI.pe._330_ ),
    .A2(\AuI.pe._341_ ),
    .B1(\AuI.pe._339_ ),
    .Y(\AuI.pe._359_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._821_  (.A(\AuI.pe._358_ ),
    .B(\AuI.pe._359_ ),
    .Y(\AuI.exponent_sub[3] ));
 sky130_fd_sc_hd__xnor2_2 \AuI.pe._822_  (.A(\AuI.operand_a[27] ),
    .B(\AuI.pe._197_ ),
    .Y(\AuI.pe._360_ ));
 sky130_fd_sc_hd__o21a_1 \AuI.pe._823_  (.A1(\AuI.pe._339_ ),
    .A2(\AuI.pe._344_ ),
    .B1(\AuI.pe._357_ ),
    .X(\AuI.pe._361_ ));
 sky130_fd_sc_hd__a31o_1 \AuI.pe._824_  (.A1(\AuI.pe._330_ ),
    .A2(\AuI.pe._341_ ),
    .A3(\AuI.pe._358_ ),
    .B1(\AuI.pe._361_ ),
    .X(\AuI.pe._362_ ));
 sky130_fd_sc_hd__xor2_1 \AuI.pe._825_  (.A(\AuI.pe._360_ ),
    .B(\AuI.pe._362_ ),
    .X(\AuI.exponent_sub[4] ));
 sky130_fd_sc_hd__a22o_1 \AuI.pe._826_  (.A1(\AuI.operand_a[27] ),
    .A2(\AuI.pe._273_ ),
    .B1(\AuI.pe._360_ ),
    .B2(\AuI.pe._362_ ),
    .X(\AuI.pe._363_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._827_  (.A1(\AuI.operand_a[27] ),
    .A2(\AuI.pe._273_ ),
    .B1(\AuI.operand_a[28] ),
    .X(\AuI.pe._364_ ));
 sky130_fd_sc_hd__a21o_1 \AuI.pe._828_  (.A1(\AuI.pe._360_ ),
    .A2(\AuI.pe._362_ ),
    .B1(\AuI.pe._364_ ),
    .X(\AuI.pe._365_ ));
 sky130_fd_sc_hd__a21bo_1 \AuI.pe._829_  (.A1(\AuI.operand_a[28] ),
    .A2(\AuI.pe._363_ ),
    .B1_N(\AuI.pe._365_ ),
    .X(\AuI.exponent_sub[5] ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._830_  (.A(\AuI.operand_a[29] ),
    .B(\AuI.pe._365_ ),
    .Y(\AuI.exponent_sub[6] ));
 sky130_fd_sc_hd__a211o_1 \AuI.pe._831_  (.A1(\AuI.pe._360_ ),
    .A2(\AuI.pe._362_ ),
    .B1(\AuI.pe._364_ ),
    .C1(\AuI.operand_a[29] ),
    .X(\AuI.pe._366_ ));
 sky130_fd_sc_hd__xnor2_1 \AuI.pe._832_  (.A(\AuI.operand_a[30] ),
    .B(\AuI.pe._366_ ),
    .Y(\AuI.exponent_sub[7] ));
 sky130_fd_sc_hd__a21o_1 \FuI._065_  (.A1(\FuI.a_operand[25] ),
    .A2(net104),
    .B1(\FuI.a_operand[26] ),
    .X(\FuI._033_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._066_  (.A1(\FuI.a_operand[28] ),
    .A2(\FuI.a_operand[29] ),
    .B1(net105),
    .X(\FuI._034_ ));
 sky130_fd_sc_hd__a31o_1 \FuI._067_  (.A1(\FuI.a_operand[27] ),
    .A2(net105),
    .A3(\FuI._033_ ),
    .B1(\FuI._034_ ),
    .X(\FuI._035_ ));
 sky130_fd_sc_hd__inv_2 \FuI._068_  (.A(\FuI.a_operand[26] ),
    .Y(\FuI._036_ ));
 sky130_fd_sc_hd__clkbuf_2 \FuI._069_  (.A(\FuI.a_operand[25] ),
    .X(\FuI._037_ ));
 sky130_fd_sc_hd__inv_2 \FuI._070_  (.A(net104),
    .Y(\FuI._038_ ));
 sky130_fd_sc_hd__and4bb_1 \FuI._071_  (.A_N(\FuI.a_operand[28] ),
    .B_N(\FuI.a_operand[29] ),
    .C(net105),
    .D(\FuI.a_operand[27] ),
    .X(\FuI._039_ ));
 sky130_fd_sc_hd__a41o_1 \FuI._072_  (.A1(\FuI._036_ ),
    .A2(\FuI._037_ ),
    .A3(\FuI._038_ ),
    .A4(\FuI._039_ ),
    .B1(\FuI._035_ ),
    .X(\FuI._040_ ));
 sky130_fd_sc_hd__o211a_1 \FuI._073_  (.A1(\FuI.a_operand[23] ),
    .A2(\FuI._035_ ),
    .B1(\FuI._040_ ),
    .C1(\FuI.a_operand[1] ),
    .X(\FuI._010_ ));
 sky130_fd_sc_hd__and2_1 \FuI._074_  (.A(\FuI.a_operand[2] ),
    .B(\FuI._040_ ),
    .X(\FuI._041_ ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._075_  (.A(\FuI._041_ ),
    .X(\FuI._014_ ));
 sky130_fd_sc_hd__a21o_1 \FuI._076_  (.A1(net104),
    .A2(\FuI.a_operand[23] ),
    .B1(\FuI.a_operand[25] ),
    .X(\FuI._042_ ));
 sky130_fd_sc_hd__and3b_1 \FuI._077_  (.A_N(\FuI._033_ ),
    .B(\FuI._039_ ),
    .C(\FuI._042_ ),
    .X(\FuI._043_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._078_  (.A1(\FuI._035_ ),
    .A2(\FuI._043_ ),
    .B1(\FuI.a_operand[3] ),
    .X(\FuI._015_ ));
 sky130_fd_sc_hd__nor2_1 \FuI._079_  (.A(\FuI.a_operand[26] ),
    .B(\FuI.a_operand[25] ),
    .Y(\FuI._044_ ));
 sky130_fd_sc_hd__and4b_1 \FuI._080_  (.A_N(\FuI.a_operand[23] ),
    .B(\FuI._044_ ),
    .C(\FuI._039_ ),
    .D(net104),
    .X(\FuI._045_ ));
 sky130_fd_sc_hd__or3_1 \FuI._081_  (.A(\FuI._035_ ),
    .B(\FuI._043_ ),
    .C(\FuI._045_ ),
    .X(\FuI._046_ ));
 sky130_fd_sc_hd__and2_1 \FuI._082_  (.A(\FuI.a_operand[4] ),
    .B(\FuI._046_ ),
    .X(\FuI._047_ ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._083_  (.A(\FuI._047_ ),
    .X(\FuI._016_ ));
 sky130_fd_sc_hd__and3_1 \FuI._084_  (.A(\FuI._038_ ),
    .B(\FuI._044_ ),
    .C(\FuI._039_ ),
    .X(\FuI._048_ ));
 sky130_fd_sc_hd__and2_1 \FuI._085_  (.A(\FuI.a_operand[23] ),
    .B(\FuI._048_ ),
    .X(\FuI._049_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._086_  (.A1(\FuI._046_ ),
    .A2(\FuI._049_ ),
    .B1(\FuI.a_operand[5] ),
    .X(\FuI._017_ ));
 sky130_fd_sc_hd__or4_1 \FuI._087_  (.A(\FuI._035_ ),
    .B(\FuI._043_ ),
    .C(\FuI._045_ ),
    .D(\FuI._048_ ),
    .X(\FuI._050_ ));
 sky130_fd_sc_hd__and2_1 \FuI._088_  (.A(\FuI.a_operand[6] ),
    .B(\FuI._050_ ),
    .X(\FuI._051_ ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._089_  (.A(\FuI._051_ ),
    .X(\FuI._018_ ));
 sky130_fd_sc_hd__buf_2 \FuI._090_  (.A(\FuI._050_ ),
    .X(\FuI._052_ ));
 sky130_fd_sc_hd__and4_1 \FuI._091_  (.A(\FuI.a_operand[26] ),
    .B(\FuI._037_ ),
    .C(net104),
    .D(\FuI.a_operand[23] ),
    .X(\FuI._053_ ));
 sky130_fd_sc_hd__o211a_1 \FuI._092_  (.A1(\FuI._052_ ),
    .A2(\FuI._053_ ),
    .B1(net105),
    .C1(\FuI.a_operand[7] ),
    .X(\FuI._019_ ));
 sky130_fd_sc_hd__or4b_2 \FuI._093_  (.A(\FuI.a_operand[27] ),
    .B(\FuI.a_operand[28] ),
    .C(\FuI.a_operand[29] ),
    .D_N(net105),
    .X(\FuI._054_ ));
 sky130_fd_sc_hd__nor2_1 \FuI._094_  (.A(\FuI._036_ ),
    .B(\FuI._054_ ),
    .Y(\FuI._055_ ));
 sky130_fd_sc_hd__clkbuf_2 \FuI._095_  (.A(\FuI._055_ ),
    .X(\FuI._056_ ));
 sky130_fd_sc_hd__and3_1 \FuI._096_  (.A(\FuI._037_ ),
    .B(net104),
    .C(\FuI._056_ ),
    .X(\FuI._057_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._097_  (.A1(\FuI._052_ ),
    .A2(\FuI._057_ ),
    .B1(\FuI.a_operand[8] ),
    .X(\FuI._020_ ));
 sky130_fd_sc_hd__or2_1 \FuI._098_  (.A(\FuI.a_operand[24] ),
    .B(\FuI.a_operand[23] ),
    .X(\FuI._058_ ));
 sky130_fd_sc_hd__and3_1 \FuI._099_  (.A(\FuI._037_ ),
    .B(\FuI._056_ ),
    .C(\FuI._058_ ),
    .X(\FuI._059_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._100_  (.A1(\FuI._052_ ),
    .A2(\FuI._059_ ),
    .B1(\FuI.a_operand[9] ),
    .X(\FuI._021_ ));
 sky130_fd_sc_hd__and2_1 \FuI._101_  (.A(\FuI._037_ ),
    .B(\FuI._055_ ),
    .X(\FuI._060_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._102_  (.A1(\FuI._052_ ),
    .A2(\FuI._060_ ),
    .B1(\FuI.a_operand[10] ),
    .X(\FuI._000_ ));
 sky130_fd_sc_hd__and2_1 \FuI._103_  (.A(net104),
    .B(\FuI.a_operand[23] ),
    .X(\FuI._061_ ));
 sky130_fd_sc_hd__and3b_1 \FuI._104_  (.A_N(\FuI._037_ ),
    .B(\FuI._061_ ),
    .C(\FuI._056_ ),
    .X(\FuI._062_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._105_  (.A1(\FuI._052_ ),
    .A2(\FuI._060_ ),
    .A3(\FuI._062_ ),
    .B1(\FuI.a_operand[11] ),
    .X(\FuI._001_ ));
 sky130_fd_sc_hd__and3b_1 \FuI._106_  (.A_N(\FuI._037_ ),
    .B(net104),
    .C(\FuI._056_ ),
    .X(\FuI._063_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._107_  (.A1(\FuI._052_ ),
    .A2(\FuI._060_ ),
    .A3(\FuI._063_ ),
    .B1(\FuI.a_operand[12] ),
    .X(\FuI._002_ ));
 sky130_fd_sc_hd__and3b_1 \FuI._108_  (.A_N(\FuI._037_ ),
    .B(\FuI._056_ ),
    .C(\FuI._058_ ),
    .X(\FuI._064_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._109_  (.A1(\FuI._052_ ),
    .A2(\FuI._060_ ),
    .A3(\FuI._064_ ),
    .B1(\FuI.a_operand[13] ),
    .X(\FuI._003_ ));
 sky130_fd_sc_hd__o21a_1 \FuI._110_  (.A1(\FuI._052_ ),
    .A2(\FuI._056_ ),
    .B1(\FuI.a_operand[14] ),
    .X(\FuI._004_ ));
 sky130_fd_sc_hd__or2b_1 \FuI._111_  (.A(\FuI.a_operand[26] ),
    .B_N(\FuI._037_ ),
    .X(\FuI._023_ ));
 sky130_fd_sc_hd__nor2_1 \FuI._112_  (.A(\FuI._023_ ),
    .B(\FuI._054_ ),
    .Y(\FuI._024_ ));
 sky130_fd_sc_hd__or3_1 \FuI._113_  (.A(\FuI._023_ ),
    .B(\FuI._061_ ),
    .C(\FuI._054_ ),
    .X(\FuI._025_ ));
 sky130_fd_sc_hd__or3_1 \FuI._114_  (.A(\FuI.a_operand[26] ),
    .B(\FuI._037_ ),
    .C(\FuI._054_ ),
    .X(\FuI._026_ ));
 sky130_fd_sc_hd__and4b_1 \FuI._115_  (.A_N(net105),
    .B(\FuI.a_operand[29] ),
    .C(\FuI.a_operand[28] ),
    .D(\FuI.a_operand[27] ),
    .X(\FuI._027_ ));
 sky130_fd_sc_hd__nand2_1 \FuI._116_  (.A(\FuI._053_ ),
    .B(\FuI._027_ ),
    .Y(\FuI._028_ ));
 sky130_fd_sc_hd__and3_1 \FuI._117_  (.A(\FuI._025_ ),
    .B(\FuI._026_ ),
    .C(\FuI._028_ ),
    .X(\FuI._029_ ));
 sky130_fd_sc_hd__o311a_1 \FuI._118_  (.A1(\FuI._050_ ),
    .A2(\FuI._056_ ),
    .A3(\FuI._024_ ),
    .B1(\FuI._029_ ),
    .C1(\FuI.a_operand[15] ),
    .X(\FuI._005_ ));
 sky130_fd_sc_hd__nand2_1 \FuI._119_  (.A(\FuI._038_ ),
    .B(\FuI._024_ ),
    .Y(\FuI._030_ ));
 sky130_fd_sc_hd__o311a_1 \FuI._120_  (.A1(\FuI._050_ ),
    .A2(\FuI._056_ ),
    .A3(\FuI._024_ ),
    .B1(\FuI._030_ ),
    .C1(\FuI.a_operand[16] ),
    .X(\FuI._006_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._121_  (.A1(\FuI._023_ ),
    .A2(\FuI._054_ ),
    .A3(\FuI._058_ ),
    .B1(\FuI.a_operand[17] ),
    .X(\FuI._031_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._122_  (.A1(\FuI._052_ ),
    .A2(\FuI._056_ ),
    .A3(\FuI._024_ ),
    .B1(\FuI._031_ ),
    .X(\FuI._007_ ));
 sky130_fd_sc_hd__o31a_1 \FuI._123_  (.A1(\FuI._052_ ),
    .A2(\FuI._056_ ),
    .A3(\FuI._024_ ),
    .B1(\FuI.a_operand[18] ),
    .X(\FuI._008_ ));
 sky130_fd_sc_hd__o211a_1 \FuI._124_  (.A1(\FuI._061_ ),
    .A2(\FuI._026_ ),
    .B1(net105),
    .C1(\FuI.a_operand[19] ),
    .X(\FuI._009_ ));
 sky130_fd_sc_hd__o211a_1 \FuI._125_  (.A1(net104),
    .A2(\FuI._026_ ),
    .B1(\FuI.a_operand[20] ),
    .C1(net105),
    .X(\FuI._011_ ));
 sky130_fd_sc_hd__o2111a_1 \FuI._126_  (.A1(\FuI._058_ ),
    .A2(\FuI._026_ ),
    .B1(\FuI._028_ ),
    .C1(\FuI.a_operand[21] ),
    .D1(net105),
    .X(\FuI._012_ ));
 sky130_fd_sc_hd__and2_1 \FuI._127_  (.A(net105),
    .B(\FuI.a_operand[22] ),
    .X(\FuI._032_ ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._128_  (.A(\FuI._032_ ),
    .X(\FuI._013_ ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._129_  (.D(\FuI._010_ ),
    .GATE_N(net135),
    .Q(\FuI.Integer[0] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._130_  (.D(\FuI._014_ ),
    .GATE_N(net136),
    .Q(\FuI.Integer[1] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._131_  (.D(\FuI._015_ ),
    .GATE_N(net137),
    .Q(\FuI.Integer[2] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._132_  (.D(\FuI._016_ ),
    .GATE_N(net138),
    .Q(\FuI.Integer[3] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._133_  (.D(\FuI._017_ ),
    .GATE_N(net139),
    .Q(\FuI.Integer[4] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._134_  (.D(\FuI._018_ ),
    .GATE_N(net140),
    .Q(\FuI.Integer[5] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._135_  (.D(\FuI._019_ ),
    .GATE_N(net141),
    .Q(\FuI.Integer[6] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._136_  (.D(\FuI._020_ ),
    .GATE_N(net142),
    .Q(\FuI.Integer[7] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._137_  (.D(\FuI._021_ ),
    .GATE_N(net143),
    .Q(\FuI.Integer[8] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._138_  (.D(\FuI._000_ ),
    .GATE_N(net144),
    .Q(\FuI.Integer[9] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._139_  (.D(\FuI._001_ ),
    .GATE_N(net145),
    .Q(\FuI.Integer[10] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._140_  (.D(\FuI._002_ ),
    .GATE_N(net146),
    .Q(\FuI.Integer[11] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._141_  (.D(\FuI._003_ ),
    .GATE_N(net147),
    .Q(\FuI.Integer[12] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._142_  (.D(\FuI._004_ ),
    .GATE_N(net148),
    .Q(\FuI.Integer[13] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._143_  (.D(\FuI._005_ ),
    .GATE_N(net149),
    .Q(\FuI.Integer[14] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._144_  (.D(\FuI._006_ ),
    .GATE_N(net150),
    .Q(\FuI.Integer[15] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._145_  (.D(\FuI._007_ ),
    .GATE_N(net151),
    .Q(\FuI.Integer[16] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._146_  (.D(\FuI._008_ ),
    .GATE_N(net152),
    .Q(\FuI.Integer[17] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._147_  (.D(\FuI._009_ ),
    .GATE_N(net153),
    .Q(\FuI.Integer[18] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._148_  (.D(\FuI._011_ ),
    .GATE_N(net154),
    .Q(\FuI.Integer[19] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._149_  (.D(\FuI._012_ ),
    .GATE_N(net155),
    .Q(\FuI.Integer[20] ));
 sky130_fd_sc_hd__dlxtn_1 \FuI._150_  (.D(\FuI._013_ ),
    .GATE_N(net156),
    .Q(\FuI.Integer[21] ));
 sky130_fd_sc_hd__conb_1 \FuI._129__135  (.LO(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__B2 (.DIODE(\AuI.Exception ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._153_  (.A(\FuI.a_operand[23] ),
    .X(\FuI.Integer[23] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._154_  (.A(net104),
    .X(\FuI.Integer[24] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._155_  (.A(\FuI.a_operand[25] ),
    .X(\FuI.Integer[25] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._156_  (.A(\FuI.a_operand[26] ),
    .X(\FuI.Integer[26] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._157_  (.A(\FuI.a_operand[27] ),
    .X(\FuI.Integer[27] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._158_  (.A(\FuI.a_operand[28] ),
    .X(\FuI.Integer[28] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._159_  (.A(\FuI.a_operand[29] ),
    .X(\FuI.Integer[29] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._160_  (.A(\FuI.a_operand[30] ),
    .X(\FuI.Integer[30] ));
 sky130_fd_sc_hd__clkbuf_1 \FuI._161_  (.A(\FuI.a_operand[31] ),
    .X(\FuI.Integer[31] ));
 sky130_fd_sc_hd__and4_1 \MuI._3423_  (.A(\MuI.b_operand[28] ),
    .B(\MuI.b_operand[27] ),
    .C(\MuI.b_operand[30] ),
    .D(\MuI.b_operand[29] ),
    .X(\MuI._0010_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3424_  (.A(\MuI.b_operand[23] ),
    .B(\MuI.b_operand[26] ),
    .C(\MuI._0010_ ),
    .X(\MuI._0021_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3425_  (.A(\MuI.a_operand[28] ),
    .B(\MuI.a_operand[27] ),
    .C(\MuI.a_operand[29] ),
    .D(\MuI.a_operand[30] ),
    .X(\MuI._0032_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3426_  (.A(\MuI.a_operand[24] ),
    .B(\MuI.a_operand[26] ),
    .C(\MuI.a_operand[25] ),
    .X(\MuI._0043_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3427_  (.A(\MuI.a_operand[23] ),
    .B(\MuI._0032_ ),
    .C(\MuI._0043_ ),
    .X(\MuI._0054_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3428_  (.A1(\MuI.b_operand[24] ),
    .A2(\MuI.b_operand[25] ),
    .A3(\MuI._0021_ ),
    .B1(\MuI._0054_ ),
    .X(\MuI._0065_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3429_  (.A(\MuI._0065_ ),
    .X(\MuI.Exception ));
 sky130_fd_sc_hd__or2_2 \MuI._3430_  (.A(\MuI.a_operand[30] ),
    .B(\MuI.b_operand[30] ),
    .X(\MuI._0086_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3431_  (.A(\MuI.a_operand[30] ),
    .B(\MuI.b_operand[30] ),
    .Y(\MuI._0097_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3432_  (.A(\MuI.a_operand[29] ),
    .B(\MuI.b_operand[29] ),
    .Y(\MuI._0108_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3433_  (.A(\MuI._0086_ ),
    .B(\MuI._0097_ ),
    .C(\MuI._0108_ ),
    .X(\MuI._0119_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3434_  (.A1(\MuI._0086_ ),
    .A2(\MuI._0097_ ),
    .B1(\MuI._0108_ ),
    .Y(\MuI._0130_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3435_  (.A(\MuI._0119_ ),
    .B(\MuI._0130_ ),
    .Y(\MuI._0141_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3436_  (.A(\MuI.a_operand[29] ),
    .B(\MuI.b_operand[29] ),
    .X(\MuI._0152_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3437_  (.A(\MuI.a_operand[28] ),
    .B(\MuI.b_operand[28] ),
    .Y(\MuI._0163_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3438_  (.A1(\MuI._0108_ ),
    .A2(\MuI._0152_ ),
    .B1_N(\MuI._0163_ ),
    .X(\MuI._0174_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3439_  (.A(\MuI.a_operand[28] ),
    .B(\MuI.b_operand[28] ),
    .X(\MuI._0185_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3440_  (.A(\MuI.a_operand[27] ),
    .B(\MuI.b_operand[27] ),
    .Y(\MuI._0196_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3441_  (.A1(\MuI._0163_ ),
    .A2(\MuI._0185_ ),
    .B1_N(\MuI._0196_ ),
    .X(\MuI._0207_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3442_  (.A(\MuI.a_operand[27] ),
    .B(\MuI.b_operand[27] ),
    .X(\MuI._0218_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3443_  (.A(\MuI.a_operand[26] ),
    .B(\MuI.b_operand[26] ),
    .Y(\MuI._0229_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3444_  (.A1(\MuI._0196_ ),
    .A2(\MuI._0218_ ),
    .B1_N(\MuI._0229_ ),
    .X(\MuI._0240_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3445_  (.A(\MuI.a_operand[26] ),
    .B(\MuI.b_operand[26] ),
    .X(\MuI._0251_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3446_  (.A(\MuI.a_operand[25] ),
    .B(\MuI.b_operand[25] ),
    .Y(\MuI._0262_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3447_  (.A1(\MuI._0229_ ),
    .A2(\MuI._0251_ ),
    .B1_N(\MuI._0262_ ),
    .X(\MuI._0273_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3448_  (.A(\MuI.a_operand[25] ),
    .B(\MuI.b_operand[25] ),
    .X(\MuI._0284_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3449_  (.A(\MuI.a_operand[24] ),
    .B(\MuI.b_operand[24] ),
    .Y(\MuI._0295_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3450_  (.A1(\MuI._0262_ ),
    .A2(\MuI._0284_ ),
    .B1_N(\MuI._0295_ ),
    .X(\MuI._0306_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3451_  (.A(\MuI.a_operand[24] ),
    .B(\MuI.b_operand[24] ),
    .X(\MuI._0317_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3452_  (.A(\MuI.a_operand[22] ),
    .X(\MuI._0328_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3453_  (.A(\MuI._0328_ ),
    .X(\MuI._0339_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3454_  (.A(\MuI._0339_ ),
    .X(\MuI._0350_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._3455_  (.A(\MuI.b_operand[22] ),
    .X(\MuI._0361_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3456_  (.A(\MuI._0361_ ),
    .X(\MuI._0372_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3457_  (.A(\MuI._0372_ ),
    .X(\MuI._0383_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3458_  (.A(\MuI._0350_ ),
    .B(\MuI._0383_ ),
    .X(\MuI._0394_ ));
 sky130_fd_sc_hd__or4_1 \MuI._3459_  (.A(\MuI.b_operand[28] ),
    .B(\MuI.b_operand[27] ),
    .C(\MuI.b_operand[30] ),
    .D(\MuI.b_operand[29] ),
    .X(\MuI._0405_ ));
 sky130_fd_sc_hd__or4_1 \MuI._3460_  (.A(\MuI.b_operand[24] ),
    .B(\MuI.b_operand[23] ),
    .C(\MuI.b_operand[26] ),
    .D(\MuI.b_operand[25] ),
    .X(\MuI._0416_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3461_  (.A(\MuI._0405_ ),
    .B(\MuI._0416_ ),
    .X(\MuI._0427_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._3462_  (.A(\MuI._0427_ ),
    .X(\MuI._0438_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3463_  (.A(\MuI._0438_ ),
    .X(\MuI._0449_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3464_  (.A(\MuI._0449_ ),
    .X(\MuI._0460_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3465_  (.A(\MuI._0460_ ),
    .X(\MuI._0471_ ));
 sky130_fd_sc_hd__nor4_4 \MuI._3466_  (.A(\MuI.a_operand[28] ),
    .B(\MuI.a_operand[27] ),
    .C(\MuI.a_operand[29] ),
    .D(\MuI.a_operand[30] ),
    .Y(\MuI._0482_ ));
 sky130_fd_sc_hd__nor4_4 \MuI._3467_  (.A(\MuI.a_operand[24] ),
    .B(\MuI.a_operand[23] ),
    .C(\MuI.a_operand[26] ),
    .D(\MuI.a_operand[25] ),
    .Y(\MuI._0493_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3468_  (.A(\MuI._0482_ ),
    .B(\MuI._0493_ ),
    .Y(\MuI._0504_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3469_  (.A(\MuI._0504_ ),
    .X(\MuI._0515_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3470_  (.A(\MuI._0515_ ),
    .X(\MuI._0526_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3471_  (.A(\MuI._0526_ ),
    .X(\MuI._0537_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3472_  (.A(\MuI._0471_ ),
    .B(\MuI._0537_ ),
    .Y(\MuI._0548_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3473_  (.A(\MuI.a_operand[21] ),
    .X(\MuI._0559_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3474_  (.A(\MuI._0559_ ),
    .X(\MuI._0570_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3475_  (.A(\MuI._0570_ ),
    .X(\MuI._0581_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3476_  (.A(\MuI._0581_ ),
    .X(\MuI._0592_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3477_  (.A(\MuI.b_operand[21] ),
    .X(\MuI._0603_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3478_  (.A(\MuI._0603_ ),
    .X(\MuI._0614_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3479_  (.A(\MuI._0614_ ),
    .X(\MuI._0625_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3480_  (.A(\MuI._0625_ ),
    .X(\MuI._0636_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3481_  (.A(\MuI._0636_ ),
    .B(\MuI._0394_ ),
    .C(\MuI._0537_ ),
    .X(\MuI._0647_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3482_  (.A1(\MuI._0636_ ),
    .A2(\MuI._0537_ ),
    .B1(\MuI._0394_ ),
    .Y(\MuI._0658_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3483_  (.A(\MuI._0647_ ),
    .B(\MuI._0658_ ),
    .Y(\MuI._0669_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3484_  (.A1(\MuI._0592_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._0669_ ),
    .B1(\MuI._0647_ ),
    .X(\MuI._0680_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3485_  (.A(\MuI._0350_ ),
    .B(\MuI._0383_ ),
    .Y(\MuI._0691_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3486_  (.A1(\MuI._0350_ ),
    .A2(\MuI._0471_ ),
    .B1(\MuI._0537_ ),
    .B2(\MuI._0383_ ),
    .X(\MuI._0702_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._3487_  (.A1(\MuI._0691_ ),
    .A2(\MuI._0548_ ),
    .B1(\MuI._0702_ ),
    .X(\MuI._0713_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3488_  (.A(\MuI._0680_ ),
    .B(\MuI._0713_ ),
    .Y(\MuI._0724_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3489_  (.A(\MuI.b_operand[19] ),
    .X(\MuI._0735_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3490_  (.A(\MuI._0735_ ),
    .X(\MuI._0746_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3491_  (.A(\MuI._0339_ ),
    .B(\MuI._0746_ ),
    .X(\MuI._0757_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3492_  (.A(\MuI.a_operand[20] ),
    .X(\MuI._0768_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3493_  (.A(\MuI._0768_ ),
    .X(\MuI._0779_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3494_  (.A(\MuI._0779_ ),
    .X(\MuI._0790_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3495_  (.A(\MuI._0790_ ),
    .X(\MuI._0801_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3496_  (.A(\MuI._0801_ ),
    .B(\MuI._0471_ ),
    .Y(\MuI._0812_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3497_  (.A1(\MuI._0350_ ),
    .A2(\MuI._0636_ ),
    .B1(\MuI._0592_ ),
    .B2(\MuI._0383_ ),
    .Y(\MuI._0823_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3498_  (.A(\MuI._0636_ ),
    .B(\MuI._0592_ ),
    .C(\MuI._0394_ ),
    .X(\MuI._0834_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3499_  (.A(\MuI._0823_ ),
    .B(\MuI._0834_ ),
    .X(\MuI._0845_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._3500_  (.A(\MuI._0812_ ),
    .B(\MuI._0845_ ),
    .X(\MuI._0856_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3501_  (.A(\MuI.b_operand[20] ),
    .X(\MuI._0867_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3502_  (.A(\MuI._0867_ ),
    .X(\MuI._0878_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3503_  (.A(\MuI._0878_ ),
    .X(\MuI._0889_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._3504_  (.A1(\MuI._0757_ ),
    .A2(\MuI._0856_ ),
    .B1(\MuI._0889_ ),
    .C1(\MuI._0537_ ),
    .X(\MuI._0900_ ));
 sky130_fd_sc_hd__inv_2 \MuI._3505_  (.A(\MuI._0900_ ),
    .Y(\MuI._0911_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._3506_  (.A1(\MuI._0812_ ),
    .A2(\MuI._0823_ ),
    .B1_N(\MuI._0834_ ),
    .X(\MuI._0922_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3507_  (.A(\MuI._0911_ ),
    .B(\MuI._0922_ ),
    .Y(\MuI._0933_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3508_  (.A(\MuI._0592_ ),
    .B(\MuI._0471_ ),
    .Y(\MuI._0944_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3509_  (.A(\MuI._0944_ ),
    .B(\MuI._0669_ ),
    .Y(\MuI._0955_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3510_  (.A(\MuI._0911_ ),
    .B(\MuI._0922_ ),
    .Y(\MuI._0966_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3511_  (.A1(\MuI._0933_ ),
    .A2(\MuI._0955_ ),
    .B1(\MuI._0966_ ),
    .Y(\MuI._0977_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3512_  (.A(\MuI._0724_ ),
    .B(\MuI._0977_ ),
    .X(\MuI._0988_ ));
 sky130_fd_sc_hd__nor3_2 \MuI._3513_  (.A(\MuI._0394_ ),
    .B(\MuI._0548_ ),
    .C(\MuI._0988_ ),
    .Y(\MuI._0999_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3514_  (.A(\MuI.a_operand[19] ),
    .X(\MuI._1010_ ));
 sky130_fd_sc_hd__buf_4 \MuI._3515_  (.A(\MuI._1010_ ),
    .X(\MuI._1021_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3516_  (.A(\MuI._1021_ ),
    .X(\MuI._1032_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3517_  (.A(\MuI._1032_ ),
    .X(\MuI._1043_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3518_  (.A1(\MuI._0636_ ),
    .A2(\MuI._0592_ ),
    .B1(\MuI._0801_ ),
    .B2(\MuI._0383_ ),
    .X(\MuI._1054_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3519_  (.A(\MuI._0383_ ),
    .B(\MuI._0636_ ),
    .C(\MuI._0592_ ),
    .D(\MuI._0801_ ),
    .X(\MuI._1065_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3520_  (.A1(\MuI._1043_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._1054_ ),
    .B1(\MuI._1065_ ),
    .X(\MuI._1076_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3521_  (.A_N(\MuI._1065_ ),
    .B(\MuI._1054_ ),
    .X(\MuI._1087_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3522_  (.A(\MuI._1043_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._1098_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3523_  (.A(\MuI._1087_ ),
    .B(\MuI._1098_ ),
    .Y(\MuI._1109_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3524_  (.A1(\MuI._0350_ ),
    .A2(\MuI._0889_ ),
    .B1(\MuI._0746_ ),
    .B2(\MuI._0526_ ),
    .Y(\MuI._1120_ ));
 sky130_fd_sc_hd__a31oi_2 \MuI._3525_  (.A1(\MuI._0889_ ),
    .A2(\MuI._0537_ ),
    .A3(\MuI._0757_ ),
    .B1(\MuI._1120_ ),
    .Y(\MuI._1131_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3526_  (.A(\MuI.b_operand[18] ),
    .X(\MuI._1142_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3527_  (.A(\MuI._1142_ ),
    .X(\MuI._1153_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3528_  (.A(\MuI._1153_ ),
    .X(\MuI._1164_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3529_  (.A(\MuI._1164_ ),
    .B(\MuI._0526_ ),
    .C(\MuI._0757_ ),
    .X(\MuI._1175_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3530_  (.A1(\MuI._1164_ ),
    .A2(\MuI._0526_ ),
    .B1(\MuI._0757_ ),
    .Y(\MuI._1186_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3531_  (.A(\MuI._1175_ ),
    .B(\MuI._1186_ ),
    .Y(\MuI._1197_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3532_  (.A(\MuI._0592_ ),
    .B(\MuI._0889_ ),
    .C(\MuI._1197_ ),
    .X(\MuI._1208_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3533_  (.A(\MuI._1175_ ),
    .B(\MuI._1208_ ),
    .X(\MuI._1219_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3534_  (.A(\MuI._1131_ ),
    .B(\MuI._1219_ ),
    .Y(\MuI._1230_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3535_  (.A(\MuI._1131_ ),
    .B(\MuI._1219_ ),
    .X(\MuI._1241_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3536_  (.A(\MuI._1230_ ),
    .B(\MuI._1241_ ),
    .X(\MuI._1252_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3537_  (.A(\MuI.b_operand[17] ),
    .X(\MuI._1263_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3538_  (.A(\MuI._1263_ ),
    .X(\MuI._1274_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3539_  (.A(\MuI._1274_ ),
    .X(\MuI._1285_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3540_  (.A(\MuI.b_operand[16] ),
    .X(\MuI._1296_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3541_  (.A(\MuI._1296_ ),
    .X(\MuI._1307_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3542_  (.A(\MuI._1307_ ),
    .X(\MuI._1318_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3543_  (.A(\MuI._0339_ ),
    .B(\MuI._1318_ ),
    .X(\MuI._1329_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3544_  (.A(\MuI._1285_ ),
    .B(\MuI._0526_ ),
    .C(\MuI._1329_ ),
    .X(\MuI._1340_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3545_  (.A1(\MuI._0592_ ),
    .A2(\MuI._0889_ ),
    .B1(\MuI._1197_ ),
    .Y(\MuI._1351_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3546_  (.A(\MuI._1208_ ),
    .B(\MuI._1351_ ),
    .X(\MuI._1362_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3547_  (.A1(\MuI._0581_ ),
    .A2(\MuI._0746_ ),
    .B1(\MuI._1164_ ),
    .B2(\MuI._0350_ ),
    .Y(\MuI._1373_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3548_  (.A(\MuI._0889_ ),
    .B(\MuI._0801_ ),
    .Y(\MuI._1384_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3549_  (.A(\MuI._0581_ ),
    .B(\MuI._1164_ ),
    .C(\MuI._0757_ ),
    .X(\MuI._1395_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._3550_  (.A1(\MuI._1373_ ),
    .A2(\MuI._1384_ ),
    .B1_N(\MuI._1395_ ),
    .X(\MuI._1406_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3551_  (.A(\MuI._1362_ ),
    .B(\MuI._1406_ ),
    .Y(\MuI._1417_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3552_  (.A1(\MuI._0636_ ),
    .A2(\MuI._0801_ ),
    .B1(\MuI._1043_ ),
    .B2(\MuI._0383_ ),
    .Y(\MuI._1428_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3553_  (.A(\MuI._0383_ ),
    .B(\MuI._0636_ ),
    .C(\MuI._0801_ ),
    .D(\MuI._1043_ ),
    .X(\MuI._1439_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3554_  (.A(\MuI._1428_ ),
    .B(\MuI._1439_ ),
    .Y(\MuI._1450_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3555_  (.A(\MuI.a_operand[18] ),
    .X(\MuI._1461_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3556_  (.A(\MuI._1461_ ),
    .X(\MuI._1472_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3557_  (.A(\MuI._1472_ ),
    .X(\MuI._1483_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3558_  (.A(\MuI._1483_ ),
    .X(\MuI._1494_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3559_  (.A(\MuI._1494_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._1505_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3560_  (.A(\MuI._1450_ ),
    .B(\MuI._1505_ ),
    .Y(\MuI._1516_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3561_  (.A(\MuI._1417_ ),
    .B(\MuI._1516_ ),
    .Y(\MuI._1527_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3562_  (.A(\MuI._1340_ ),
    .B(\MuI._1527_ ),
    .Y(\MuI._1538_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3563_  (.A(\MuI._1109_ ),
    .B(\MuI._1252_ ),
    .Y(\MuI._1549_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3564_  (.A(\MuI._1538_ ),
    .B(\MuI._1549_ ),
    .Y(\MuI._1560_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3565_  (.A(\MuI._1230_ ),
    .B(\MuI._1560_ ),
    .Y(\MuI._1571_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3566_  (.A1(\MuI._1109_ ),
    .A2(\MuI._1252_ ),
    .B1(\MuI._1571_ ),
    .Y(\MuI._1582_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3567_  (.A(\MuI._1076_ ),
    .B(\MuI._1582_ ),
    .Y(\MuI._1593_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._3568_  (.A_N(\MuI._0757_ ),
    .B(\MuI._0889_ ),
    .C(\MuI._0537_ ),
    .Y(\MuI._1604_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._3569_  (.A(\MuI._0856_ ),
    .B(\MuI._1604_ ),
    .Y(\MuI._1615_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3570_  (.A(\MuI._0966_ ),
    .B_N(\MuI._0933_ ),
    .X(\MuI._1626_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3571_  (.A(\MuI._1626_ ),
    .B(\MuI._0955_ ),
    .Y(\MuI._1637_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3572_  (.A(\MuI._1593_ ),
    .B(\MuI._1615_ ),
    .C(\MuI._1637_ ),
    .Y(\MuI._1648_ ));
 sky130_fd_sc_hd__inv_2 \MuI._3573_  (.A(\MuI._1076_ ),
    .Y(\MuI._1659_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3574_  (.A(\MuI._1659_ ),
    .B(\MuI._1582_ ),
    .Y(\MuI._1670_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3575_  (.A1(\MuI._1131_ ),
    .A2(\MuI._1219_ ),
    .A3(\MuI._1560_ ),
    .B1(\MuI._1670_ ),
    .X(\MuI._1681_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3576_  (.A1(\MuI._1593_ ),
    .A2(\MuI._1615_ ),
    .B1(\MuI._1637_ ),
    .X(\MuI._1692_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3577_  (.A(\MuI._1648_ ),
    .B(\MuI._1692_ ),
    .X(\MuI._1703_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3578_  (.A(\MuI._1681_ ),
    .B(\MuI._1703_ ),
    .Y(\MuI._1714_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3579_  (.A(\MuI._0724_ ),
    .B(\MuI._0977_ ),
    .Y(\MuI._1725_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3580_  (.A(\MuI._0988_ ),
    .B(\MuI._1725_ ),
    .Y(\MuI._1736_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3581_  (.A1(\MuI._1648_ ),
    .A2(\MuI._1714_ ),
    .B1(\MuI._1736_ ),
    .Y(\MuI._1747_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3582_  (.A(\MuI._1681_ ),
    .B(\MuI._1703_ ),
    .Y(\MuI._1758_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3583_  (.A(\MuI._1340_ ),
    .B(\MuI._1527_ ),
    .X(\MuI._1769_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3584_  (.A(\MuI._1538_ ),
    .B(\MuI._1769_ ),
    .Y(\MuI._1780_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3585_  (.A(\MuI.b_operand[15] ),
    .X(\MuI._1791_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3586_  (.A(\MuI._1791_ ),
    .X(\MuI._1802_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3587_  (.A(\MuI._1802_ ),
    .X(\MuI._1813_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3588_  (.A(\MuI._1813_ ),
    .B(\MuI._0515_ ),
    .C(\MuI._1329_ ),
    .X(\MuI._1824_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3589_  (.A1(\MuI._1813_ ),
    .A2(\MuI._0515_ ),
    .B1(\MuI._1329_ ),
    .Y(\MuI._1835_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3590_  (.A(\MuI._1824_ ),
    .B(\MuI._1835_ ),
    .Y(\MuI._1846_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3591_  (.A1(\MuI._0592_ ),
    .A2(\MuI._1285_ ),
    .A3(\MuI._1846_ ),
    .B1(\MuI._1824_ ),
    .X(\MuI._1857_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3592_  (.A1(\MuI._0350_ ),
    .A2(\MuI._1285_ ),
    .B1(\MuI._1318_ ),
    .B2(\MuI._0526_ ),
    .Y(\MuI._1868_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3593_  (.A(\MuI._1340_ ),
    .B(\MuI._1868_ ),
    .Y(\MuI._1879_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._3594_  (.A_N(\MuI._1329_ ),
    .B(\MuI._1285_ ),
    .C(\MuI._0537_ ),
    .X(\MuI._1890_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3595_  (.A(\MuI._1857_ ),
    .B(\MuI._1879_ ),
    .Y(\MuI._1901_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3596_  (.A(\MuI._1901_ ),
    .B(\MuI._1890_ ),
    .X(\MuI._1912_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3597_  (.A(\MuI._0581_ ),
    .B(\MuI._0746_ ),
    .C(\MuI._0801_ ),
    .D(\MuI._1153_ ),
    .X(\MuI._1923_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3598_  (.A1(\MuI._0746_ ),
    .A2(\MuI._0801_ ),
    .B1(\MuI._1164_ ),
    .B2(\MuI._0581_ ),
    .Y(\MuI._1934_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3599_  (.A(\MuI._1923_ ),
    .B(\MuI._1934_ ),
    .Y(\MuI._1945_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3600_  (.A(\MuI._0889_ ),
    .B(\MuI._1043_ ),
    .C(\MuI._1945_ ),
    .X(\MuI._1956_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3601_  (.A(\MuI._1395_ ),
    .B(\MuI._1373_ ),
    .Y(\MuI._1967_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3602_  (.A(\MuI._1967_ ),
    .B(\MuI._1384_ ),
    .Y(\MuI._1978_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._3603_  (.A1(\MuI._1923_ ),
    .A2(\MuI._1956_ ),
    .B1(\MuI._1978_ ),
    .X(\MuI._1989_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3604_  (.A(\MuI._1978_ ),
    .B(\MuI._1923_ ),
    .C(\MuI._1956_ ),
    .X(\MuI._2000_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3605_  (.A_N(\MuI._1989_ ),
    .B(\MuI._2000_ ),
    .X(\MuI._2011_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3606_  (.A1(\MuI._0636_ ),
    .A2(\MuI._1043_ ),
    .B1(\MuI._1494_ ),
    .B2(\MuI._0383_ ),
    .Y(\MuI._2022_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3607_  (.A(\MuI._0383_ ),
    .B(\MuI._0625_ ),
    .C(\MuI._1043_ ),
    .D(\MuI._1494_ ),
    .X(\MuI._2033_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3608_  (.A(\MuI._2022_ ),
    .B(\MuI._2033_ ),
    .X(\MuI._2044_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3609_  (.A(\MuI.a_operand[17] ),
    .X(\MuI._2055_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3610_  (.A(\MuI._2055_ ),
    .X(\MuI._2066_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3611_  (.A(\MuI._2066_ ),
    .X(\MuI._2077_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3612_  (.A(\MuI._2077_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._2088_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3613_  (.A(\MuI._2044_ ),
    .B(\MuI._2088_ ),
    .X(\MuI._2099_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3614_  (.A(\MuI._2011_ ),
    .B(\MuI._2099_ ),
    .Y(\MuI._2110_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3615_  (.A(\MuI._1912_ ),
    .B(\MuI._2110_ ),
    .Y(\MuI._2121_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3616_  (.A1(\MuI._1857_ ),
    .A2(\MuI._1879_ ),
    .A3(\MuI._1890_ ),
    .B1(\MuI._2121_ ),
    .X(\MuI._2132_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3617_  (.A_N(\MuI._1780_ ),
    .B(\MuI._2132_ ),
    .X(\MuI._2143_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3618_  (.A(\MuI._1417_ ),
    .B_N(\MuI._1516_ ),
    .X(\MuI._2154_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._3619_  (.A1(\MuI._1362_ ),
    .A2(\MuI._1406_ ),
    .B1(\MuI._2154_ ),
    .X(\MuI._2165_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3620_  (.A(\MuI._2143_ ),
    .B(\MuI._2165_ ),
    .Y(\MuI._2176_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3621_  (.A1(\MuI._1494_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._1450_ ),
    .B1(\MuI._1439_ ),
    .X(\MuI._2187_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._3622_  (.A(\MuI._1780_ ),
    .B(\MuI._2165_ ),
    .C_N(\MuI._2132_ ),
    .X(\MuI._2198_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3623_  (.A1(\MuI._2176_ ),
    .A2(\MuI._2187_ ),
    .B1_N(\MuI._2198_ ),
    .X(\MuI._2209_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3624_  (.A(\MuI._1593_ ),
    .B(\MuI._1615_ ),
    .X(\MuI._2220_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3625_  (.A(\MuI._2176_ ),
    .B(\MuI._2187_ ),
    .X(\MuI._2231_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3626_  (.A(\MuI._1538_ ),
    .B(\MuI._1549_ ),
    .X(\MuI._2242_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3627_  (.A(\MuI._1560_ ),
    .B(\MuI._2242_ ),
    .Y(\MuI._2253_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3628_  (.A(\MuI._2231_ ),
    .B(\MuI._2253_ ),
    .X(\MuI._2264_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3629_  (.A(\MuI._2220_ ),
    .B(\MuI._2264_ ),
    .X(\MuI._2275_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3630_  (.A(\MuI._2220_ ),
    .B(\MuI._2264_ ),
    .X(\MuI._2286_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3631_  (.A1(\MuI._2209_ ),
    .A2(\MuI._2275_ ),
    .B1(\MuI._2286_ ),
    .Y(\MuI._2297_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3632_  (.A(\MuI._1758_ ),
    .B(\MuI._2297_ ),
    .Y(\MuI._2308_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3633_  (.A(\MuI.a_operand[6] ),
    .X(\MuI._2319_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3634_  (.A(\MuI._2319_ ),
    .X(\MuI._2330_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3635_  (.A(\MuI.a_operand[8] ),
    .X(\MuI._2341_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3636_  (.A(\MuI._2341_ ),
    .X(\MuI._2352_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3637_  (.A(\MuI._2352_ ),
    .X(\MuI._2363_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3638_  (.A(\MuI.a_operand[7] ),
    .X(\MuI._2374_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3639_  (.A(\MuI._2374_ ),
    .X(\MuI._2385_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3640_  (.A1(\MuI.b_operand[21] ),
    .A2(\MuI._2363_ ),
    .B1(\MuI._2385_ ),
    .B2(\MuI.b_operand[22] ),
    .X(\MuI._2396_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3641_  (.A(\MuI.b_operand[22] ),
    .B(\MuI.b_operand[21] ),
    .C(\MuI._2363_ ),
    .X(\MuI._2407_ ));
 sky130_fd_sc_hd__a32o_1 \MuI._3642_  (.A1(\MuI._2330_ ),
    .A2(\MuI._0460_ ),
    .A3(\MuI._2396_ ),
    .B1(\MuI._2407_ ),
    .B2(\MuI._2385_ ),
    .X(\MuI._2418_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3643_  (.A(\MuI.a_operand[13] ),
    .X(\MuI._2429_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3644_  (.A(\MuI._2429_ ),
    .X(\MuI._2440_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3645_  (.A(\MuI.a_operand[12] ),
    .X(\MuI._2451_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3646_  (.A(\MuI._1307_ ),
    .B(\MuI._1802_ ),
    .C(\MuI._2440_ ),
    .D(\MuI._2451_ ),
    .X(\MuI._2462_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3647_  (.A(\MuI.b_operand[17] ),
    .X(\MuI._2473_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3648_  (.A(\MuI.a_operand[11] ),
    .X(\MuI._2484_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3649_  (.A(\MuI._2484_ ),
    .X(\MuI._2495_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3650_  (.A(\MuI._2473_ ),
    .B(\MuI._2495_ ),
    .Y(\MuI._2506_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3651_  (.A(\MuI._1791_ ),
    .X(\MuI._2517_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3652_  (.A(\MuI._2429_ ),
    .X(\MuI._2528_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3653_  (.A(\MuI._2451_ ),
    .X(\MuI._2539_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3654_  (.A(\MuI._1296_ ),
    .X(\MuI._2550_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3655_  (.A1(\MuI._2517_ ),
    .A2(\MuI._2528_ ),
    .B1(\MuI._2539_ ),
    .B2(\MuI._2550_ ),
    .Y(\MuI._2561_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3656_  (.A(\MuI._2462_ ),
    .B(\MuI._2506_ ),
    .C(\MuI._2561_ ),
    .X(\MuI._2572_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3657_  (.A(\MuI.b_operand[14] ),
    .X(\MuI._2583_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3658_  (.A(\MuI._2528_ ),
    .X(\MuI._2594_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3659_  (.A(\MuI.a_operand[15] ),
    .X(\MuI._2605_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3660_  (.A(\MuI._2605_ ),
    .X(\MuI._2616_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3661_  (.A(\MuI._2616_ ),
    .X(\MuI._2627_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3662_  (.A(\MuI.b_operand[12] ),
    .X(\MuI._2638_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3663_  (.A(\MuI._2638_ ),
    .X(\MuI._2649_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3664_  (.A(\MuI.a_operand[14] ),
    .X(\MuI._2660_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3665_  (.A(\MuI._2660_ ),
    .X(\MuI._2671_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3666_  (.A(\MuI._2671_ ),
    .X(\MuI._2682_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3667_  (.A(\MuI.b_operand[13] ),
    .X(\MuI._2693_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3668_  (.A(\MuI._2693_ ),
    .X(\MuI._2704_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3669_  (.A1(\MuI._2627_ ),
    .A2(\MuI._2649_ ),
    .B1(\MuI._2682_ ),
    .B2(\MuI._2704_ ),
    .X(\MuI._2715_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3670_  (.A(\MuI._2704_ ),
    .B(\MuI._2616_ ),
    .C(\MuI._2649_ ),
    .D(\MuI._2671_ ),
    .X(\MuI._2726_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3671_  (.A1(\MuI._2583_ ),
    .A2(\MuI._2594_ ),
    .A3(\MuI._2715_ ),
    .B1(\MuI._2726_ ),
    .X(\MuI._2736_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3672_  (.A1(\MuI._2462_ ),
    .A2(\MuI._2561_ ),
    .B1(\MuI._2506_ ),
    .Y(\MuI._2743_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3673_  (.A(\MuI._2572_ ),
    .B(\MuI._2736_ ),
    .C(\MuI._2743_ ),
    .Y(\MuI._2748_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3674_  (.A(\MuI.b_operand[15] ),
    .X(\MuI._2754_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3675_  (.A(\MuI._1307_ ),
    .B(\MuI._2754_ ),
    .C(\MuI._2451_ ),
    .D(\MuI._2484_ ),
    .X(\MuI._2759_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3676_  (.A(\MuI.a_operand[10] ),
    .X(\MuI._2765_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3677_  (.A(\MuI._2765_ ),
    .X(\MuI._2773_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3678_  (.A(\MuI._1263_ ),
    .B(\MuI._2773_ ),
    .Y(\MuI._2778_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3679_  (.A1(\MuI._2517_ ),
    .A2(\MuI._2539_ ),
    .B1(\MuI._2495_ ),
    .B2(\MuI._2550_ ),
    .Y(\MuI._2779_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3680_  (.A(\MuI._2759_ ),
    .B(\MuI._2778_ ),
    .C(\MuI._2779_ ),
    .X(\MuI._2780_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3681_  (.A(\MuI._2759_ ),
    .B_N(\MuI._2780_ ),
    .X(\MuI._2781_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3682_  (.A1(\MuI._2572_ ),
    .A2(\MuI._2743_ ),
    .B1(\MuI._2736_ ),
    .X(\MuI._2782_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3683_  (.A(\MuI._2748_ ),
    .B(\MuI._2781_ ),
    .C(\MuI._2782_ ),
    .Y(\MuI._2783_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3684_  (.A1(\MuI._2748_ ),
    .A2(\MuI._2782_ ),
    .B1(\MuI._2781_ ),
    .X(\MuI._2784_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3685_  (.A(\MuI.a_operand[9] ),
    .X(\MuI._2785_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3686_  (.A(\MuI._2785_ ),
    .X(\MuI._2786_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3687_  (.A(\MuI._2786_ ),
    .X(\MuI._2787_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3688_  (.A(\MuI._2550_ ),
    .B(\MuI._2517_ ),
    .C(\MuI._2495_ ),
    .D(\MuI._2773_ ),
    .X(\MuI._2788_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3689_  (.A(\MuI._2484_ ),
    .X(\MuI._2789_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3690_  (.A(\MuI.a_operand[10] ),
    .X(\MuI._2790_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3691_  (.A(\MuI._2790_ ),
    .X(\MuI._2791_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3692_  (.A1(\MuI._2517_ ),
    .A2(\MuI._2789_ ),
    .B1(\MuI._2791_ ),
    .B2(\MuI._1318_ ),
    .Y(\MuI._2792_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3693_  (.A(\MuI._2788_ ),
    .B(\MuI._2792_ ),
    .Y(\MuI._2793_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3694_  (.A1(\MuI._1274_ ),
    .A2(\MuI._2787_ ),
    .A3(\MuI._2793_ ),
    .B1(\MuI._2788_ ),
    .X(\MuI._2794_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3695_  (.A1(\MuI._2759_ ),
    .A2(\MuI._2779_ ),
    .B1(\MuI._2778_ ),
    .Y(\MuI._2795_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3696_  (.A(\MuI.b_operand[14] ),
    .X(\MuI._2796_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3697_  (.A(\MuI._2539_ ),
    .X(\MuI._2797_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3698_  (.A(\MuI._2796_ ),
    .B(\MuI._2797_ ),
    .Y(\MuI._2798_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3699_  (.A(\MuI.b_operand[13] ),
    .X(\MuI._2799_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3700_  (.A(\MuI._2799_ ),
    .X(\MuI._2800_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3701_  (.A1(\MuI._2649_ ),
    .A2(\MuI._2682_ ),
    .B1(\MuI._2528_ ),
    .B2(\MuI._2800_ ),
    .Y(\MuI._2801_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3702_  (.A(\MuI._2693_ ),
    .X(\MuI._2802_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3703_  (.A(\MuI._2638_ ),
    .X(\MuI._2803_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3704_  (.A(\MuI._2802_ ),
    .B(\MuI._2803_ ),
    .C(\MuI._2671_ ),
    .D(\MuI._2528_ ),
    .X(\MuI._2804_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._3705_  (.A1(\MuI._2798_ ),
    .A2(\MuI._2801_ ),
    .B1_N(\MuI._2804_ ),
    .Y(\MuI._2805_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3706_  (.A1(\MuI._2780_ ),
    .A2(\MuI._2795_ ),
    .B1(\MuI._2805_ ),
    .X(\MuI._2806_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3707_  (.A(\MuI._2780_ ),
    .B(\MuI._2805_ ),
    .C(\MuI._2795_ ),
    .Y(\MuI._2807_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3708_  (.A1(\MuI._2794_ ),
    .A2(\MuI._2806_ ),
    .B1_N(\MuI._2807_ ),
    .X(\MuI._2808_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3709_  (.A(\MuI._2783_ ),
    .B(\MuI._2784_ ),
    .C(\MuI._2808_ ),
    .X(\MuI._2809_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3710_  (.A1(\MuI._2783_ ),
    .A2(\MuI._2784_ ),
    .B1(\MuI._2808_ ),
    .Y(\MuI._2810_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._3711_  (.A(\MuI.b_operand[18] ),
    .X(\MuI._2811_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3712_  (.A(\MuI.b_operand[19] ),
    .B(\MuI._2811_ ),
    .C(\MuI._2773_ ),
    .D(\MuI._2786_ ),
    .X(\MuI._2812_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3713_  (.A(\MuI._2811_ ),
    .X(\MuI._2813_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3714_  (.A(\MuI.b_operand[19] ),
    .X(\MuI._2814_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3715_  (.A1(\MuI._2813_ ),
    .A2(\MuI._2773_ ),
    .B1(\MuI._2786_ ),
    .B2(\MuI._2814_ ),
    .Y(\MuI._2815_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._3716_  (.A_N(\MuI._2812_ ),
    .B_N(\MuI._2815_ ),
    .C(\MuI._0867_ ),
    .D(\MuI._2363_ ),
    .X(\MuI._2816_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3717_  (.A(\MuI.b_operand[20] ),
    .X(\MuI._2817_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._3718_  (.A1_N(\MuI._2817_ ),
    .A2_N(\MuI._2363_ ),
    .B1(\MuI._2812_ ),
    .B2(\MuI._2815_ ),
    .X(\MuI._2818_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3719_  (.A(\MuI._2816_ ),
    .B(\MuI._2818_ ),
    .Y(\MuI._2819_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3720_  (.A(\MuI._2814_ ),
    .B(\MuI._1142_ ),
    .C(\MuI._2786_ ),
    .D(\MuI._2352_ ),
    .X(\MuI._2820_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3721_  (.A1(\MuI._2813_ ),
    .A2(\MuI._2786_ ),
    .B1(\MuI._2363_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._2821_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._3722_  (.A_N(\MuI._2820_ ),
    .B_N(\MuI._2821_ ),
    .C(\MuI._0867_ ),
    .D(\MuI._2385_ ),
    .X(\MuI._2822_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3723_  (.A(\MuI._2820_ ),
    .B(\MuI._2822_ ),
    .Y(\MuI._2823_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3724_  (.A(\MuI._2819_ ),
    .B(\MuI._2823_ ),
    .Y(\MuI._2824_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3725_  (.A1(\MuI._0614_ ),
    .A2(\MuI._2385_ ),
    .B1(\MuI._2330_ ),
    .B2(\MuI._0361_ ),
    .Y(\MuI._2825_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3726_  (.A(\MuI.b_operand[22] ),
    .X(\MuI._2826_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3727_  (.A(\MuI._2826_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._2385_ ),
    .D(\MuI._2330_ ),
    .X(\MuI._2827_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3728_  (.A(\MuI._2825_ ),
    .B(\MuI._2827_ ),
    .Y(\MuI._2828_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3729_  (.A(\MuI.a_operand[5] ),
    .X(\MuI._2829_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3730_  (.A(\MuI._2829_ ),
    .X(\MuI._2830_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3731_  (.A(\MuI._2830_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._2831_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3732_  (.A(\MuI._2828_ ),
    .B(\MuI._2831_ ),
    .Y(\MuI._2832_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3733_  (.A(\MuI._2824_ ),
    .B(\MuI._2832_ ),
    .Y(\MuI._2833_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3734_  (.A(\MuI._2809_ ),
    .B(\MuI._2810_ ),
    .C(\MuI._2833_ ),
    .X(\MuI._2834_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3735_  (.A(\MuI._2809_ ),
    .B_N(\MuI._2834_ ),
    .X(\MuI._2835_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3736_  (.A(\MuI.b_operand[10] ),
    .X(\MuI._2836_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3737_  (.A(\MuI.b_operand[9] ),
    .X(\MuI._2837_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3738_  (.A(\MuI._2837_ ),
    .X(\MuI._2838_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3739_  (.A(\MuI._1461_ ),
    .B(\MuI._2055_ ),
    .C(\MuI._2836_ ),
    .D(\MuI._2838_ ),
    .X(\MuI._2839_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3740_  (.A(\MuI.a_operand[16] ),
    .X(\MuI._2840_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3741_  (.A(\MuI.b_operand[11] ),
    .X(\MuI._2841_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3742_  (.A(\MuI._2840_ ),
    .B(\MuI._2841_ ),
    .Y(\MuI._2842_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3743_  (.A(\MuI._2055_ ),
    .X(\MuI._2843_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3744_  (.A(\MuI.b_operand[10] ),
    .X(\MuI._2844_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3745_  (.A(\MuI._2837_ ),
    .X(\MuI._2845_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3746_  (.A1(\MuI._2843_ ),
    .A2(\MuI._2844_ ),
    .B1(\MuI._2845_ ),
    .B2(\MuI._1472_ ),
    .Y(\MuI._2846_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3747_  (.A(\MuI._2839_ ),
    .B(\MuI._2842_ ),
    .C(\MuI._2846_ ),
    .X(\MuI._2847_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3748_  (.A1(\MuI._2839_ ),
    .A2(\MuI._2846_ ),
    .B1(\MuI._2842_ ),
    .Y(\MuI._2848_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3749_  (.A(\MuI._2627_ ),
    .X(\MuI._2849_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3750_  (.A(\MuI.b_operand[11] ),
    .X(\MuI._2850_ ));
 sky130_fd_sc_hd__buf_4 \MuI._3751_  (.A(\MuI._2850_ ),
    .X(\MuI._2851_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3752_  (.A(\MuI.a_operand[16] ),
    .X(\MuI._2852_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3753_  (.A(\MuI.b_operand[10] ),
    .X(\MuI._2853_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3754_  (.A(\MuI.b_operand[9] ),
    .X(\MuI._2854_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3755_  (.A1(\MuI._2852_ ),
    .A2(\MuI._2853_ ),
    .B1(\MuI._2854_ ),
    .B2(\MuI._2055_ ),
    .X(\MuI._2855_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3756_  (.A(\MuI._2055_ ),
    .B(\MuI._2852_ ),
    .C(\MuI.b_operand[10] ),
    .D(\MuI._2837_ ),
    .X(\MuI._2856_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3757_  (.A1(\MuI._2849_ ),
    .A2(\MuI._2851_ ),
    .A3(\MuI._2855_ ),
    .B1(\MuI._2856_ ),
    .X(\MuI._2857_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3758_  (.A(\MuI._2847_ ),
    .B(\MuI._2848_ ),
    .C(\MuI._2857_ ),
    .Y(\MuI._2858_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3759_  (.A1(\MuI._2847_ ),
    .A2(\MuI._2848_ ),
    .B1(\MuI._2857_ ),
    .X(\MuI._2859_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3760_  (.A(\MuI._2796_ ),
    .X(\MuI._2860_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3761_  (.A(\MuI._2860_ ),
    .B(\MuI._2594_ ),
    .Y(\MuI._2861_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3762_  (.A_N(\MuI._2726_ ),
    .B(\MuI._2715_ ),
    .X(\MuI._2862_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3763_  (.A(\MuI._2861_ ),
    .B(\MuI._2862_ ),
    .Y(\MuI._2863_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3764_  (.A(\MuI._2858_ ),
    .B(\MuI._2859_ ),
    .C(\MuI._2863_ ),
    .Y(\MuI._2864_ ));
 sky130_fd_sc_hd__nand2_2 \MuI._3765_  (.A(\MuI._2858_ ),
    .B(\MuI._2864_ ),
    .Y(\MuI._2865_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3766_  (.A(\MuI.b_operand[7] ),
    .X(\MuI._2866_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3767_  (.A(\MuI._2866_ ),
    .X(\MuI._2867_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3768_  (.A(\MuI.b_operand[6] ),
    .X(\MuI._2868_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3769_  (.A(\MuI._2868_ ),
    .X(\MuI._2869_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3770_  (.A(\MuI._0779_ ),
    .B(\MuI._1021_ ),
    .C(\MuI._2867_ ),
    .D(\MuI._2869_ ),
    .X(\MuI._2870_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3771_  (.A(\MuI.b_operand[8] ),
    .X(\MuI._2871_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3772_  (.A(\MuI._1483_ ),
    .B(\MuI._2871_ ),
    .Y(\MuI._2872_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3773_  (.A(\MuI._2866_ ),
    .X(\MuI._2873_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3774_  (.A(\MuI._2873_ ),
    .X(\MuI._2874_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3775_  (.A(\MuI._2868_ ),
    .X(\MuI._2875_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3776_  (.A(\MuI._2875_ ),
    .X(\MuI._2876_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3777_  (.A1(\MuI._1021_ ),
    .A2(\MuI._2874_ ),
    .B1(\MuI._2876_ ),
    .B2(\MuI._0790_ ),
    .Y(\MuI._2877_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3778_  (.A(\MuI._2870_ ),
    .B(\MuI._2872_ ),
    .C(\MuI._2877_ ),
    .X(\MuI._2878_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3779_  (.A(\MuI._2870_ ),
    .B_N(\MuI._2878_ ),
    .X(\MuI._2879_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3780_  (.A(\MuI.b_operand[3] ),
    .X(\MuI._2880_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3781_  (.A(\MuI._2880_ ),
    .X(\MuI._2881_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3782_  (.A(\MuI._2881_ ),
    .X(\MuI._2882_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3783_  (.A(\MuI._0328_ ),
    .B(\MuI._2882_ ),
    .Y(\MuI._2883_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3784_  (.A(\MuI.b_operand[4] ),
    .X(\MuI._2884_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3785_  (.A(\MuI._2884_ ),
    .X(\MuI._2885_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3786_  (.A(\MuI._2885_ ),
    .X(\MuI._2886_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3787_  (.A1(\MuI._0482_ ),
    .A2(\MuI._0493_ ),
    .B1_N(\MuI._2886_ ),
    .X(\MuI._2887_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3788_  (.A(\MuI._2883_ ),
    .B(\MuI._2887_ ),
    .Y(\MuI._2888_ ));
 sky130_fd_sc_hd__or4_4 \MuI._3789_  (.A(\MuI.a_operand[28] ),
    .B(\MuI.a_operand[27] ),
    .C(\MuI.a_operand[29] ),
    .D(\MuI.a_operand[30] ),
    .X(\MuI._2889_ ));
 sky130_fd_sc_hd__or3_4 \MuI._3790_  (.A(\MuI.a_operand[24] ),
    .B(\MuI.a_operand[23] ),
    .C(\MuI.a_operand[26] ),
    .X(\MuI._2890_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._3791_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._2882_ ),
    .X(\MuI._2891_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3792_  (.A(\MuI._2884_ ),
    .X(\MuI._2892_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3793_  (.A(\MuI._0328_ ),
    .B(\MuI._2892_ ),
    .X(\MuI._2893_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3794_  (.A(\MuI._0559_ ),
    .X(\MuI._2894_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3795_  (.A(\MuI.b_operand[5] ),
    .X(\MuI._2895_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3796_  (.A(\MuI._2894_ ),
    .B(\MuI._2895_ ),
    .X(\MuI._2896_ ));
 sky130_fd_sc_hd__o221a_1 \MuI._3797_  (.A1(\MuI._2883_ ),
    .A2(\MuI._2887_ ),
    .B1(\MuI._2891_ ),
    .B2(\MuI._2893_ ),
    .C1(\MuI._2896_ ),
    .X(\MuI._2897_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3798_  (.A(\MuI._2871_ ),
    .X(\MuI._2898_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3799_  (.A(\MuI._1032_ ),
    .B(\MuI._2898_ ),
    .Y(\MuI._2899_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3800_  (.A(\MuI._2894_ ),
    .B(\MuI._0768_ ),
    .C(\MuI._2867_ ),
    .D(\MuI._2869_ ),
    .X(\MuI._2900_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3801_  (.A1(\MuI._0779_ ),
    .A2(\MuI._2874_ ),
    .B1(\MuI._2876_ ),
    .B2(\MuI._2894_ ),
    .Y(\MuI._2901_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3802_  (.A(\MuI._2900_ ),
    .B(\MuI._2901_ ),
    .Y(\MuI._2902_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3803_  (.A(\MuI._2899_ ),
    .B(\MuI._2902_ ),
    .Y(\MuI._2903_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3804_  (.A(\MuI._2888_ ),
    .B(\MuI._2897_ ),
    .C(\MuI._2903_ ),
    .X(\MuI._2904_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3805_  (.A1(\MuI._2888_ ),
    .A2(\MuI._2897_ ),
    .B1(\MuI._2903_ ),
    .Y(\MuI._2905_ ));
 sky130_fd_sc_hd__a21boi_2 \MuI._3806_  (.A1(\MuI._2879_ ),
    .A2(\MuI._2904_ ),
    .B1_N(\MuI._2905_ ),
    .Y(\MuI._2906_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3807_  (.A(\MuI._2066_ ),
    .B(\MuI._2850_ ),
    .Y(\MuI._2907_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3808_  (.A(\MuI._1010_ ),
    .B(\MuI._1472_ ),
    .C(\MuI._2836_ ),
    .D(\MuI._2838_ ),
    .X(\MuI._2908_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3809_  (.A1(\MuI._1472_ ),
    .A2(\MuI._2844_ ),
    .B1(\MuI._2845_ ),
    .B2(\MuI._1010_ ),
    .X(\MuI._2909_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3810_  (.A_N(\MuI._2908_ ),
    .B(\MuI._2909_ ),
    .X(\MuI._2910_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._3811_  (.A(\MuI._2907_ ),
    .B(\MuI._2910_ ),
    .Y(\MuI._2911_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3812_  (.A(\MuI._2839_ ),
    .B_N(\MuI._2847_ ),
    .X(\MuI._2912_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._3813_  (.A(\MuI._2911_ ),
    .B(\MuI._2912_ ),
    .X(\MuI._2913_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3814_  (.A(\MuI._2682_ ),
    .X(\MuI._2914_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3815_  (.A(\MuI._2860_ ),
    .B(\MuI._2914_ ),
    .Y(\MuI._2915_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3816_  (.A(\MuI._2840_ ),
    .X(\MuI._2916_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3817_  (.A(\MuI._2916_ ),
    .B(\MuI._2704_ ),
    .C(\MuI._2627_ ),
    .D(\MuI._2649_ ),
    .X(\MuI._2917_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3818_  (.A(\MuI.b_operand[12] ),
    .X(\MuI._2918_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3819_  (.A(\MuI._2918_ ),
    .X(\MuI._2919_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3820_  (.A1(\MuI._2704_ ),
    .A2(\MuI._2627_ ),
    .B1(\MuI._2919_ ),
    .B2(\MuI._2916_ ),
    .X(\MuI._2920_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3821_  (.A_N(\MuI._2917_ ),
    .B(\MuI._2920_ ),
    .X(\MuI._2921_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._3822_  (.A(\MuI._2915_ ),
    .B(\MuI._2921_ ),
    .Y(\MuI._2922_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._3823_  (.A(\MuI._2913_ ),
    .B(\MuI._2922_ ),
    .X(\MuI._2923_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._3824_  (.A(\MuI._2906_ ),
    .B(\MuI._2923_ ),
    .Y(\MuI._2924_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3825_  (.A_N(\MuI._2906_ ),
    .B(\MuI._2923_ ),
    .X(\MuI._2925_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._3826_  (.A1(\MuI._2865_ ),
    .A2(\MuI._2924_ ),
    .B1(\MuI._2925_ ),
    .Y(\MuI._2926_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3827_  (.A(\MuI._2462_ ),
    .B_N(\MuI._2572_ ),
    .X(\MuI._2927_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3828_  (.A1(\MuI._2860_ ),
    .A2(\MuI._2914_ ),
    .A3(\MuI._2920_ ),
    .B1(\MuI._2917_ ),
    .X(\MuI._2928_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3829_  (.A(\MuI._1274_ ),
    .B(\MuI._2797_ ),
    .Y(\MuI._2929_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3830_  (.A(\MuI._1307_ ),
    .B(\MuI._1802_ ),
    .C(\MuI._2440_ ),
    .X(\MuI._2930_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3831_  (.A1(\MuI._1802_ ),
    .A2(\MuI._2671_ ),
    .B1(\MuI._2440_ ),
    .B2(\MuI._1307_ ),
    .X(\MuI._2931_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3832_  (.A1(\MuI._2682_ ),
    .A2(\MuI._2930_ ),
    .B1_N(\MuI._2931_ ),
    .X(\MuI._2932_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3833_  (.A(\MuI._2929_ ),
    .B(\MuI._2932_ ),
    .X(\MuI._2933_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3834_  (.A(\MuI._2928_ ),
    .B(\MuI._2933_ ),
    .X(\MuI._2934_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3835_  (.A(\MuI._2927_ ),
    .B(\MuI._2934_ ),
    .Y(\MuI._2935_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3836_  (.A(\MuI._2748_ ),
    .B(\MuI._2783_ ),
    .X(\MuI._2936_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3837_  (.A(\MuI._2935_ ),
    .B(\MuI._2936_ ),
    .Y(\MuI._2937_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3838_  (.A(\MuI.b_operand[19] ),
    .B(\MuI._2811_ ),
    .C(\MuI._2484_ ),
    .D(\MuI._2773_ ),
    .X(\MuI._2938_ ));
 sky130_fd_sc_hd__buf_2 \MuI._3839_  (.A(\MuI.b_operand[19] ),
    .X(\MuI._2939_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3840_  (.A1(\MuI._1142_ ),
    .A2(\MuI._2495_ ),
    .B1(\MuI._2791_ ),
    .B2(\MuI._2939_ ),
    .Y(\MuI._2940_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3841_  (.A(\MuI._2938_ ),
    .B(\MuI._2940_ ),
    .Y(\MuI._2941_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3842_  (.A(\MuI._0867_ ),
    .B(\MuI._2787_ ),
    .Y(\MuI._2942_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3843_  (.A(\MuI._2941_ ),
    .B(\MuI._2942_ ),
    .Y(\MuI._2943_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3844_  (.A(\MuI._2812_ ),
    .B(\MuI._2816_ ),
    .Y(\MuI._2944_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3845_  (.A(\MuI._2943_ ),
    .B(\MuI._2944_ ),
    .Y(\MuI._2945_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3846_  (.A1(\MuI._2385_ ),
    .A2(\MuI._2407_ ),
    .B1_N(\MuI._2396_ ),
    .X(\MuI._2946_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3847_  (.A(\MuI._2330_ ),
    .B(\MuI._0438_ ),
    .Y(\MuI._2947_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3848_  (.A(\MuI._2946_ ),
    .B(\MuI._2947_ ),
    .X(\MuI._2948_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3849_  (.A(\MuI._2945_ ),
    .B(\MuI._2948_ ),
    .X(\MuI._2949_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3850_  (.A(\MuI._2945_ ),
    .B(\MuI._2948_ ),
    .Y(\MuI._2950_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3851_  (.A(\MuI._2949_ ),
    .B(\MuI._2950_ ),
    .X(\MuI._2951_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3852_  (.A(\MuI._2937_ ),
    .B(\MuI._2951_ ),
    .Y(\MuI._2952_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3853_  (.A(\MuI._2926_ ),
    .B(\MuI._2952_ ),
    .X(\MuI._2953_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3854_  (.A(\MuI._2926_ ),
    .B(\MuI._2952_ ),
    .Y(\MuI._2954_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3855_  (.A1(\MuI._2835_ ),
    .A2(\MuI._2953_ ),
    .B1(\MuI._2954_ ),
    .X(\MuI._2955_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3856_  (.A_N(\MuI._2944_ ),
    .B(\MuI._2943_ ),
    .X(\MuI._2956_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3857_  (.A(\MuI._2956_ ),
    .B(\MuI._2949_ ),
    .Y(\MuI._2957_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3858_  (.A(\MuI._2955_ ),
    .B(\MuI._2957_ ),
    .Y(\MuI._2958_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3859_  (.A1(\MuI._2956_ ),
    .A2(\MuI._2949_ ),
    .B1(\MuI._2955_ ),
    .Y(\MuI._2959_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3860_  (.A1(\MuI._2418_ ),
    .A2(\MuI._2958_ ),
    .B1_N(\MuI._2959_ ),
    .X(\MuI._2960_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3861_  (.A(\MuI._0779_ ),
    .B(\MuI._2871_ ),
    .Y(\MuI._2961_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._3862_  (.A(\MuI._0328_ ),
    .B(\MuI._2894_ ),
    .C(\MuI._2874_ ),
    .D(\MuI._2869_ ),
    .Y(\MuI._2962_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3863_  (.A1(\MuI._2894_ ),
    .A2(\MuI._2867_ ),
    .B1(\MuI._2869_ ),
    .B2(\MuI._0328_ ),
    .X(\MuI._2963_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._3864_  (.A_N(\MuI._2961_ ),
    .B(\MuI._2962_ ),
    .C(\MuI._2963_ ),
    .Y(\MuI._2964_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3865_  (.A1(\MuI._2962_ ),
    .A2(\MuI._2963_ ),
    .B1_N(\MuI._2961_ ),
    .X(\MuI._2965_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3866_  (.A(\MuI.b_operand[5] ),
    .X(\MuI._2966_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3867_  (.A(\MuI._2966_ ),
    .X(\MuI._2967_ ));
 sky130_fd_sc_hd__o311a_1 \MuI._3868_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._2893_ ),
    .C1(\MuI._2967_ ),
    .X(\MuI._2968_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3869_  (.A1(\MuI._2964_ ),
    .A2(\MuI._2965_ ),
    .B1(\MuI._2968_ ),
    .X(\MuI._2969_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3870_  (.A1(\MuI._1032_ ),
    .A2(\MuI._2898_ ),
    .A3(\MuI._2902_ ),
    .B1(\MuI._2900_ ),
    .X(\MuI._2970_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3871_  (.A(\MuI._2968_ ),
    .B(\MuI._2964_ ),
    .C(\MuI._2965_ ),
    .Y(\MuI._2971_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3872_  (.A1(\MuI._2969_ ),
    .A2(\MuI._2970_ ),
    .B1_N(\MuI._2971_ ),
    .X(\MuI._2972_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3873_  (.A(\MuI._1472_ ),
    .B(\MuI._2841_ ),
    .Y(\MuI._2973_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3874_  (.A(\MuI._0768_ ),
    .B(\MuI._1010_ ),
    .C(\MuI._2844_ ),
    .D(\MuI._2838_ ),
    .X(\MuI._2974_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3875_  (.A(\MuI._2853_ ),
    .X(\MuI._2975_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3876_  (.A(\MuI._2838_ ),
    .X(\MuI._2976_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._3877_  (.A1(\MuI._1010_ ),
    .A2(\MuI._2975_ ),
    .B1(\MuI._2976_ ),
    .B2(\MuI._0779_ ),
    .Y(\MuI._2977_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3878_  (.A(\MuI._2973_ ),
    .B(\MuI._2974_ ),
    .C(\MuI._2977_ ),
    .X(\MuI._2978_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3879_  (.A1(\MuI._2974_ ),
    .A2(\MuI._2977_ ),
    .B1(\MuI._2973_ ),
    .Y(\MuI._2979_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3880_  (.A1(\MuI._2066_ ),
    .A2(\MuI._2850_ ),
    .A3(\MuI._2909_ ),
    .B1(\MuI._2908_ ),
    .X(\MuI._2980_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3881_  (.A(\MuI._2978_ ),
    .B(\MuI._2979_ ),
    .C(\MuI._2980_ ),
    .Y(\MuI._2981_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3882_  (.A1(\MuI._2978_ ),
    .A2(\MuI._2979_ ),
    .B1(\MuI._2980_ ),
    .X(\MuI._2982_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3883_  (.A(\MuI.b_operand[14] ),
    .B(\MuI._2616_ ),
    .Y(\MuI._2983_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3884_  (.A(\MuI._2843_ ),
    .B(\MuI._2840_ ),
    .C(\MuI._2799_ ),
    .D(\MuI._2918_ ),
    .X(\MuI._2984_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3885_  (.A1(\MuI._2840_ ),
    .A2(\MuI._2802_ ),
    .B1(\MuI._2649_ ),
    .B2(\MuI._2843_ ),
    .Y(\MuI._2985_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3886_  (.A(\MuI._2984_ ),
    .B(\MuI._2985_ ),
    .Y(\MuI._2986_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3887_  (.A(\MuI._2983_ ),
    .B(\MuI._2986_ ),
    .Y(\MuI._2987_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3888_  (.A(\MuI._2981_ ),
    .B(\MuI._2982_ ),
    .C(\MuI._2987_ ),
    .Y(\MuI._2988_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3889_  (.A1(\MuI._2981_ ),
    .A2(\MuI._2982_ ),
    .B1(\MuI._2987_ ),
    .X(\MuI._2989_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3890_  (.A(\MuI._2911_ ),
    .B(\MuI._2912_ ),
    .X(\MuI._2990_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3891_  (.A(\MuI._2913_ ),
    .B(\MuI._2922_ ),
    .X(\MuI._2991_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3892_  (.A(\MuI._2972_ ),
    .B(\MuI._2988_ ),
    .C(\MuI._2989_ ),
    .Y(\MuI._2992_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3893_  (.A1(\MuI._2988_ ),
    .A2(\MuI._2989_ ),
    .B1(\MuI._2972_ ),
    .X(\MuI._2993_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._3894_  (.A1(\MuI._2990_ ),
    .A2(\MuI._2991_ ),
    .B1(\MuI._2992_ ),
    .C1(\MuI._2993_ ),
    .X(\MuI._2994_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3895_  (.A1(\MuI._2972_ ),
    .A2(\MuI._2988_ ),
    .A3(\MuI._2989_ ),
    .B1(\MuI._2994_ ),
    .X(\MuI._2995_ ));
 sky130_fd_sc_hd__a32o_1 \MuI._3896_  (.A1(\MuI._1274_ ),
    .A2(\MuI._2797_ ),
    .A3(\MuI._2931_ ),
    .B1(\MuI._2930_ ),
    .B2(\MuI._2914_ ),
    .X(\MuI._2996_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._3897_  (.A1(\MuI._2983_ ),
    .A2(\MuI._2985_ ),
    .B1_N(\MuI._2984_ ),
    .Y(\MuI._2997_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3898_  (.A(\MuI._1263_ ),
    .B(\MuI._2528_ ),
    .Y(\MuI._2998_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._3899_  (.A(\MuI._1307_ ),
    .B(\MuI._1802_ ),
    .C(\MuI._2616_ ),
    .D(\MuI._2671_ ),
    .Y(\MuI._2999_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._3900_  (.A(\MuI.b_operand[16] ),
    .X(\MuI._3000_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3901_  (.A1(\MuI._2754_ ),
    .A2(\MuI._2605_ ),
    .B1(\MuI._2660_ ),
    .B2(\MuI._3000_ ),
    .X(\MuI._3001_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._3902_  (.A_N(\MuI._2998_ ),
    .B(\MuI._2999_ ),
    .C(\MuI._3001_ ),
    .Y(\MuI._3002_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3903_  (.A1(\MuI._2999_ ),
    .A2(\MuI._3001_ ),
    .B1_N(\MuI._2998_ ),
    .X(\MuI._3003_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3904_  (.A(\MuI._2997_ ),
    .B(\MuI._3002_ ),
    .C(\MuI._3003_ ),
    .Y(\MuI._3004_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3905_  (.A1(\MuI._3002_ ),
    .A2(\MuI._3003_ ),
    .B1(\MuI._2997_ ),
    .X(\MuI._3005_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3906_  (.A(\MuI._2996_ ),
    .B(\MuI._3004_ ),
    .C(\MuI._3005_ ),
    .X(\MuI._3006_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3907_  (.A1(\MuI._3004_ ),
    .A2(\MuI._3005_ ),
    .B1(\MuI._2996_ ),
    .Y(\MuI._3007_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3908_  (.A(\MuI._3006_ ),
    .B(\MuI._3007_ ),
    .X(\MuI._3008_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3909_  (.A(\MuI._2928_ ),
    .B(\MuI._2933_ ),
    .X(\MuI._3009_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3910_  (.A1(\MuI._2927_ ),
    .A2(\MuI._2934_ ),
    .B1(\MuI._3009_ ),
    .Y(\MuI._3010_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3911_  (.A(\MuI._3008_ ),
    .B(\MuI._3010_ ),
    .Y(\MuI._3011_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3912_  (.A(\MuI._2817_ ),
    .B(\MuI._2787_ ),
    .C(\MuI._2941_ ),
    .X(\MuI._3012_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3913_  (.A(\MuI._2939_ ),
    .B(\MuI._2811_ ),
    .C(\MuI._2451_ ),
    .D(\MuI._2495_ ),
    .X(\MuI._3013_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3914_  (.A1(\MuI._2813_ ),
    .A2(\MuI._2539_ ),
    .B1(\MuI._2495_ ),
    .B2(\MuI._2814_ ),
    .Y(\MuI._3014_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3915_  (.A(\MuI._3013_ ),
    .B(\MuI._3014_ ),
    .Y(\MuI._3015_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3916_  (.A(\MuI._0867_ ),
    .B(\MuI._2791_ ),
    .Y(\MuI._3016_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3917_  (.A(\MuI._3015_ ),
    .B(\MuI._3016_ ),
    .Y(\MuI._3017_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3918_  (.A1(\MuI._2938_ ),
    .A2(\MuI._3012_ ),
    .B1(\MuI._3017_ ),
    .Y(\MuI._3018_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3919_  (.A(\MuI._2938_ ),
    .B(\MuI._3012_ ),
    .C(\MuI._3017_ ),
    .X(\MuI._3019_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3920_  (.A(\MuI._3018_ ),
    .B(\MuI._3019_ ),
    .Y(\MuI._3020_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3921_  (.A1(\MuI._0603_ ),
    .A2(\MuI._2787_ ),
    .B1(\MuI._2363_ ),
    .B2(\MuI._2826_ ),
    .X(\MuI._3021_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3922_  (.A1(\MuI._2787_ ),
    .A2(\MuI._2407_ ),
    .B1_N(\MuI._3021_ ),
    .X(\MuI._3022_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3923_  (.A(\MuI._2385_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._3023_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3924_  (.A(\MuI._3022_ ),
    .B(\MuI._3023_ ),
    .Y(\MuI._3024_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3925_  (.A(\MuI._3020_ ),
    .B(\MuI._3024_ ),
    .X(\MuI._3025_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3926_  (.A(\MuI._3011_ ),
    .B(\MuI._3025_ ),
    .Y(\MuI._3026_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3927_  (.A(\MuI._2995_ ),
    .B(\MuI._3026_ ),
    .X(\MuI._3027_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3928_  (.A(\MuI._2995_ ),
    .B(\MuI._3026_ ),
    .Y(\MuI._3028_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3929_  (.A(\MuI._2935_ ),
    .B(\MuI._2936_ ),
    .X(\MuI._3029_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._3930_  (.A1(\MuI._2937_ ),
    .A2(\MuI._2951_ ),
    .B1(\MuI._3029_ ),
    .Y(\MuI._3030_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3931_  (.A_N(\MuI._3028_ ),
    .B(\MuI._3030_ ),
    .X(\MuI._3031_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._3932_  (.A1(\MuI._3020_ ),
    .A2(\MuI._3024_ ),
    .B1(\MuI._3018_ ),
    .X(\MuI._3032_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._3933_  (.A1(\MuI._3027_ ),
    .A2(\MuI._3031_ ),
    .B1_N(\MuI._3032_ ),
    .X(\MuI._3033_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._3934_  (.A(\MuI._3027_ ),
    .B(\MuI._3031_ ),
    .C_N(\MuI._3032_ ),
    .X(\MuI._3034_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3935_  (.A_N(\MuI._3033_ ),
    .B(\MuI._3034_ ),
    .X(\MuI._3035_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._3936_  (.A1_N(\MuI._2787_ ),
    .A2_N(\MuI._2407_ ),
    .B1(\MuI._3022_ ),
    .B2(\MuI._3023_ ),
    .X(\MuI._3036_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3937_  (.A(\MuI._3035_ ),
    .B(\MuI._3036_ ),
    .Y(\MuI._3037_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3938_  (.A(\MuI._2962_ ),
    .B(\MuI._2964_ ),
    .Y(\MuI._3038_ ));
 sky130_fd_sc_hd__inv_2 \MuI._3939_  (.A(\MuI._3038_ ),
    .Y(\MuI._3039_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3940_  (.A(\MuI._1010_ ),
    .B(\MuI.b_operand[11] ),
    .Y(\MuI._3040_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3941_  (.A(\MuI._0559_ ),
    .B(\MuI._0768_ ),
    .C(\MuI._2853_ ),
    .D(\MuI._2854_ ),
    .X(\MuI._3041_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._3942_  (.A1(\MuI._0768_ ),
    .A2(\MuI._2836_ ),
    .B1(\MuI._2845_ ),
    .B2(\MuI._0559_ ),
    .Y(\MuI._3042_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3943_  (.A(\MuI._3040_ ),
    .B(\MuI._3041_ ),
    .C(\MuI._3042_ ),
    .X(\MuI._3043_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._3944_  (.A1(\MuI._3041_ ),
    .A2(\MuI._3042_ ),
    .B1(\MuI._3040_ ),
    .Y(\MuI._3044_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._3945_  (.A1(\MuI._2973_ ),
    .A2(\MuI._2977_ ),
    .B1_N(\MuI._2974_ ),
    .Y(\MuI._3045_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3946_  (.A(\MuI._3043_ ),
    .B(\MuI._3044_ ),
    .C(\MuI._3045_ ),
    .Y(\MuI._3046_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3947_  (.A1(\MuI._3043_ ),
    .A2(\MuI._3044_ ),
    .B1(\MuI._3045_ ),
    .X(\MuI._3047_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3948_  (.A(\MuI._2916_ ),
    .B(\MuI._2796_ ),
    .Y(\MuI._3048_ ));
 sky130_fd_sc_hd__and4_1 \MuI._3949_  (.A(\MuI._1461_ ),
    .B(\MuI._2055_ ),
    .C(\MuI._2693_ ),
    .D(\MuI._2638_ ),
    .X(\MuI._3049_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3950_  (.A1(\MuI._2055_ ),
    .A2(\MuI._2693_ ),
    .B1(\MuI._2918_ ),
    .B2(\MuI._1472_ ),
    .X(\MuI._3050_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._3951_  (.A_N(\MuI._3049_ ),
    .B(\MuI._3050_ ),
    .X(\MuI._3051_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3952_  (.A(\MuI._3048_ ),
    .B(\MuI._3051_ ),
    .Y(\MuI._3052_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3953_  (.A(\MuI._3046_ ),
    .B(\MuI._3047_ ),
    .C(\MuI._3052_ ),
    .X(\MuI._3053_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._3954_  (.A1(\MuI._3046_ ),
    .A2(\MuI._3047_ ),
    .B1(\MuI._3052_ ),
    .Y(\MuI._3054_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3955_  (.A(\MuI._0581_ ),
    .B(\MuI._2898_ ),
    .Y(\MuI._3055_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3956_  (.A(\MuI._0328_ ),
    .B(\MuI._2874_ ),
    .X(\MuI._3056_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._3957_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._2876_ ),
    .X(\MuI._3057_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3958_  (.A(\MuI._3056_ ),
    .B(\MuI._3057_ ),
    .X(\MuI._3058_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3959_  (.A(\MuI._3055_ ),
    .B(\MuI._3058_ ),
    .Y(\MuI._3059_ ));
 sky130_fd_sc_hd__or4b_1 \MuI._3960_  (.A(\MuI._3039_ ),
    .B(\MuI._3053_ ),
    .C(\MuI._3054_ ),
    .D_N(\MuI._3059_ ),
    .X(\MuI._3060_ ));
 sky130_fd_sc_hd__a2bb2o_1 \MuI._3961_  (.A1_N(\MuI._3053_ ),
    .A2_N(\MuI._3054_ ),
    .B1(\MuI._3038_ ),
    .B2(\MuI._3059_ ),
    .X(\MuI._3061_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3962_  (.A(\MuI._3060_ ),
    .B(\MuI._3061_ ),
    .X(\MuI._3062_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3963_  (.A(\MuI._2981_ ),
    .B(\MuI._2988_ ),
    .Y(\MuI._3063_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._3964_  (.A(\MuI._3062_ ),
    .B(\MuI._3063_ ),
    .X(\MuI._3064_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3965_  (.A(\MuI._3056_ ),
    .B(\MuI._3057_ ),
    .X(\MuI._3065_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3966_  (.A1(\MuI._0581_ ),
    .A2(\MuI._2898_ ),
    .A3(\MuI._3058_ ),
    .B1(\MuI._3065_ ),
    .X(\MuI._3066_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3967_  (.A(\MuI._2898_ ),
    .B(\MuI._0515_ ),
    .C(\MuI._3056_ ),
    .X(\MuI._3067_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._3968_  (.A1(\MuI._0350_ ),
    .A2(\MuI._2898_ ),
    .B1(\MuI._2874_ ),
    .B2(\MuI._0515_ ),
    .Y(\MuI._3068_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._3969_  (.A(\MuI._3067_ ),
    .B(\MuI._3068_ ),
    .Y(\MuI._3069_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3970_  (.A(\MuI._3066_ ),
    .B(\MuI._3069_ ),
    .Y(\MuI._3070_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3971_  (.A(\MuI._3064_ ),
    .B(\MuI._3070_ ),
    .Y(\MuI._3071_ ));
 sky130_fd_sc_hd__and2_1 \MuI._3972_  (.A(\MuI._2967_ ),
    .B(\MuI._0515_ ),
    .X(\MuI._3072_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3973_  (.A(\MuI._2971_ ),
    .B(\MuI._2969_ ),
    .C(\MuI._2970_ ),
    .Y(\MuI._3073_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3974_  (.A1(\MuI._2971_ ),
    .A2(\MuI._2969_ ),
    .B1(\MuI._2970_ ),
    .X(\MuI._3074_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3975_  (.A(\MuI._3072_ ),
    .B(\MuI._3073_ ),
    .C(\MuI._3074_ ),
    .X(\MuI._3075_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3976_  (.A(\MuI._3039_ ),
    .B(\MuI._3059_ ),
    .Y(\MuI._3076_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._3977_  (.A1(\MuI._2992_ ),
    .A2(\MuI._2993_ ),
    .B1(\MuI._2990_ ),
    .C1(\MuI._2991_ ),
    .Y(\MuI._3077_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3978_  (.A(\MuI._3075_ ),
    .B(\MuI._3076_ ),
    .Y(\MuI._3078_ ));
 sky130_fd_sc_hd__or3_1 \MuI._3979_  (.A(\MuI._2994_ ),
    .B(\MuI._3077_ ),
    .C(\MuI._3078_ ),
    .X(\MuI._3079_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3980_  (.A1(\MuI._3075_ ),
    .A2(\MuI._3076_ ),
    .B1_N(\MuI._3079_ ),
    .X(\MuI._3080_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3981_  (.A(\MuI._3071_ ),
    .B(\MuI._3080_ ),
    .Y(\MuI._3081_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._3982_  (.A(\MuI._3028_ ),
    .B(\MuI._3030_ ),
    .X(\MuI._3082_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._3983_  (.A(\MuI._3071_ ),
    .B(\MuI._3080_ ),
    .Y(\MuI._3083_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3984_  (.A(\MuI._3082_ ),
    .B(\MuI._3083_ ),
    .X(\MuI._3084_ ));
 sky130_fd_sc_hd__or2_1 \MuI._3985_  (.A(\MuI._3008_ ),
    .B(\MuI._3010_ ),
    .X(\MuI._3085_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._3986_  (.A(\MuI._3011_ ),
    .B_N(\MuI._3025_ ),
    .X(\MuI._3086_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3987_  (.A(\MuI._3046_ ),
    .B(\MuI._3047_ ),
    .C(\MuI._3052_ ),
    .Y(\MuI._3087_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._3988_  (.A_N(\MuI._3039_ ),
    .B_N(\MuI._3054_ ),
    .C(\MuI._3059_ ),
    .D(\MuI._3087_ ),
    .X(\MuI._3088_ ));
 sky130_fd_sc_hd__and3_1 \MuI._3989_  (.A(\MuI._3060_ ),
    .B(\MuI._3061_ ),
    .C(\MuI._3063_ ),
    .X(\MuI._3089_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3990_  (.A(\MuI._2999_ ),
    .B(\MuI._3002_ ),
    .Y(\MuI._3090_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._3991_  (.A(\MuI._2916_ ),
    .X(\MuI._3091_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._3992_  (.A1(\MuI._3091_ ),
    .A2(\MuI._2860_ ),
    .A3(\MuI._3050_ ),
    .B1(\MuI._3049_ ),
    .X(\MuI._3092_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._3993_  (.A(\MuI._2473_ ),
    .B(\MuI._2682_ ),
    .Y(\MuI._3093_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._3994_  (.A(\MuI._1318_ ),
    .B(\MuI._1813_ ),
    .C(\MuI._2916_ ),
    .D(\MuI._2627_ ),
    .Y(\MuI._3094_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._3995_  (.A1(\MuI._2517_ ),
    .A2(\MuI._2916_ ),
    .B1(\MuI._2627_ ),
    .B2(\MuI._1318_ ),
    .X(\MuI._3095_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._3996_  (.A_N(\MuI._3093_ ),
    .B(\MuI._3094_ ),
    .C(\MuI._3095_ ),
    .Y(\MuI._3096_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._3997_  (.A1(\MuI._3094_ ),
    .A2(\MuI._3095_ ),
    .B1_N(\MuI._3093_ ),
    .X(\MuI._3097_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._3998_  (.A(\MuI._3092_ ),
    .B(\MuI._3096_ ),
    .C(\MuI._3097_ ),
    .Y(\MuI._3098_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._3999_  (.A1(\MuI._3096_ ),
    .A2(\MuI._3097_ ),
    .B1(\MuI._3092_ ),
    .X(\MuI._3099_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4000_  (.A(\MuI._3090_ ),
    .B(\MuI._3098_ ),
    .C(\MuI._3099_ ),
    .Y(\MuI._3100_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4001_  (.A1(\MuI._3098_ ),
    .A2(\MuI._3099_ ),
    .B1(\MuI._3090_ ),
    .X(\MuI._3101_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4002_  (.A1(\MuI._2996_ ),
    .A2(\MuI._3005_ ),
    .B1_N(\MuI._3004_ ),
    .X(\MuI._3102_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4003_  (.A(\MuI._3100_ ),
    .B(\MuI._3101_ ),
    .C(\MuI._3102_ ),
    .X(\MuI._3103_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4004_  (.A1(\MuI._3100_ ),
    .A2(\MuI._3101_ ),
    .B1(\MuI._3102_ ),
    .Y(\MuI._3104_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4005_  (.A(\MuI._2814_ ),
    .B(\MuI._1142_ ),
    .C(\MuI._2528_ ),
    .D(\MuI._2539_ ),
    .X(\MuI._3105_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4006_  (.A1(\MuI._1153_ ),
    .A2(\MuI._2528_ ),
    .B1(\MuI._2797_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._3106_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4007_  (.A(\MuI._3105_ ),
    .B(\MuI._3106_ ),
    .Y(\MuI._3107_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4008_  (.A(\MuI._2817_ ),
    .B(\MuI._2789_ ),
    .Y(\MuI._3108_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4009_  (.A(\MuI._3107_ ),
    .B(\MuI._3108_ ),
    .Y(\MuI._3109_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4010_  (.A1(\MuI._3014_ ),
    .A2(\MuI._3016_ ),
    .B1_N(\MuI._3013_ ),
    .X(\MuI._3110_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4011_  (.A(\MuI._3109_ ),
    .B(\MuI._3110_ ),
    .Y(\MuI._3111_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4012_  (.A1(\MuI.b_operand[21] ),
    .A2(\MuI._2791_ ),
    .B1(\MuI._2787_ ),
    .B2(\MuI.b_operand[22] ),
    .X(\MuI._3112_ ));
 sky130_fd_sc_hd__inv_2 \MuI._4013_  (.A(\MuI._3112_ ),
    .Y(\MuI._3113_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4014_  (.A(\MuI._0361_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._2791_ ),
    .D(\MuI._2787_ ),
    .X(\MuI._3114_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4015_  (.A(\MuI._3113_ ),
    .B(\MuI._3114_ ),
    .Y(\MuI._3115_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4016_  (.A(\MuI._2363_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._3116_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4017_  (.A(\MuI._3115_ ),
    .B(\MuI._3116_ ),
    .Y(\MuI._3117_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4018_  (.A(\MuI._3111_ ),
    .B(\MuI._3117_ ),
    .Y(\MuI._3118_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4019_  (.A(\MuI._3103_ ),
    .B(\MuI._3104_ ),
    .C(\MuI._3118_ ),
    .X(\MuI._3119_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4020_  (.A1(\MuI._3103_ ),
    .A2(\MuI._3104_ ),
    .B1(\MuI._3118_ ),
    .Y(\MuI._3120_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._4021_  (.A1(\MuI._3088_ ),
    .A2(\MuI._3089_ ),
    .B1(\MuI._3119_ ),
    .C1(\MuI._3120_ ),
    .X(\MuI._3121_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._4022_  (.A1(\MuI._3119_ ),
    .A2(\MuI._3120_ ),
    .B1(\MuI._3088_ ),
    .C1(\MuI._3089_ ),
    .Y(\MuI._3122_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._4023_  (.A1(\MuI._3085_ ),
    .A2(\MuI._3086_ ),
    .B1(\MuI._3121_ ),
    .C1(\MuI._3122_ ),
    .Y(\MuI._3123_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._4024_  (.A1(\MuI._3121_ ),
    .A2(\MuI._3122_ ),
    .B1(\MuI._3085_ ),
    .C1(\MuI._3086_ ),
    .X(\MuI._3124_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4025_  (.A(\MuI._3123_ ),
    .B(\MuI._3124_ ),
    .Y(\MuI._3125_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4026_  (.A(\MuI._2898_ ),
    .B(\MuI._0526_ ),
    .Y(\MuI._3126_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._4027_  (.A1(\MuI._3040_ ),
    .A2(\MuI._3042_ ),
    .B1_N(\MuI._3041_ ),
    .Y(\MuI._3127_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4028_  (.A(\MuI._0790_ ),
    .B(\MuI._2851_ ),
    .Y(\MuI._3128_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._4029_  (.A(\MuI._0339_ ),
    .B(\MuI._0570_ ),
    .C(\MuI._2975_ ),
    .D(\MuI._2976_ ),
    .Y(\MuI._3129_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4030_  (.A1(\MuI._0570_ ),
    .A2(\MuI._2975_ ),
    .B1(\MuI._2976_ ),
    .B2(\MuI._0339_ ),
    .X(\MuI._3130_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._4031_  (.A_N(\MuI._3128_ ),
    .B(\MuI._3129_ ),
    .C(\MuI._3130_ ),
    .Y(\MuI._3131_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4032_  (.A1(\MuI._3129_ ),
    .A2(\MuI._3130_ ),
    .B1_N(\MuI._3128_ ),
    .X(\MuI._3132_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4033_  (.A(\MuI._3127_ ),
    .B(\MuI._3131_ ),
    .C(\MuI._3132_ ),
    .Y(\MuI._3133_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4034_  (.A1(\MuI._3131_ ),
    .A2(\MuI._3132_ ),
    .B1(\MuI._3127_ ),
    .X(\MuI._3134_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4035_  (.A(\MuI._2077_ ),
    .B(\MuI._2583_ ),
    .Y(\MuI._3135_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4036_  (.A(\MuI._1032_ ),
    .B(\MuI._1483_ ),
    .C(\MuI._2800_ ),
    .D(\MuI._2919_ ),
    .X(\MuI._3136_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4037_  (.A1(\MuI._1494_ ),
    .A2(\MuI._2800_ ),
    .B1(\MuI._2919_ ),
    .B2(\MuI._1032_ ),
    .Y(\MuI._3137_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4038_  (.A(\MuI._3136_ ),
    .B(\MuI._3137_ ),
    .Y(\MuI._3138_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4039_  (.A(\MuI._3135_ ),
    .B(\MuI._3138_ ),
    .Y(\MuI._3139_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4040_  (.A(\MuI._3133_ ),
    .B(\MuI._3134_ ),
    .C(\MuI._3139_ ),
    .Y(\MuI._3140_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4041_  (.A1(\MuI._3133_ ),
    .A2(\MuI._3134_ ),
    .B1(\MuI._3139_ ),
    .X(\MuI._3141_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._4042_  (.A(\MuI._3066_ ),
    .B(\MuI._3069_ ),
    .C(\MuI._3140_ ),
    .D(\MuI._3141_ ),
    .Y(\MuI._3142_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4043_  (.A1(\MuI._3066_ ),
    .A2(\MuI._3069_ ),
    .B1(\MuI._3140_ ),
    .B2(\MuI._3141_ ),
    .X(\MuI._3143_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4044_  (.A(\MuI._3046_ ),
    .B(\MuI._3087_ ),
    .Y(\MuI._3144_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4045_  (.A(\MuI._3142_ ),
    .B(\MuI._3143_ ),
    .C(\MuI._3144_ ),
    .Y(\MuI._3145_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4046_  (.A1(\MuI._3142_ ),
    .A2(\MuI._3143_ ),
    .B1(\MuI._3144_ ),
    .X(\MuI._3146_ ));
 sky130_fd_sc_hd__or4bb_1 \MuI._4047_  (.A(\MuI._3056_ ),
    .B(\MuI._3126_ ),
    .C_N(\MuI._3145_ ),
    .D_N(\MuI._3146_ ),
    .X(\MuI._3147_ ));
 sky130_fd_sc_hd__a2bb2o_1 \MuI._4048_  (.A1_N(\MuI._3056_ ),
    .A2_N(\MuI._3126_ ),
    .B1(\MuI._3145_ ),
    .B2(\MuI._3146_ ),
    .X(\MuI._3148_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4049_  (.A(\MuI._3147_ ),
    .B(\MuI._3148_ ),
    .Y(\MuI._3149_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4050_  (.A(\MuI._3062_ ),
    .B(\MuI._3063_ ),
    .Y(\MuI._3150_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4051_  (.A(\MuI._3089_ ),
    .B(\MuI._3150_ ),
    .C(\MuI._3070_ ),
    .X(\MuI._3151_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4052_  (.A(\MuI._3149_ ),
    .B(\MuI._3151_ ),
    .X(\MuI._3152_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4053_  (.A(\MuI._3125_ ),
    .B(\MuI._3152_ ),
    .Y(\MuI._3153_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4054_  (.A1(\MuI._3081_ ),
    .A2(\MuI._3084_ ),
    .B1(\MuI._3153_ ),
    .Y(\MuI._3154_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4055_  (.A(\MuI._3153_ ),
    .B(\MuI._3081_ ),
    .C(\MuI._3084_ ),
    .X(\MuI._3155_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4056_  (.A(\MuI._3154_ ),
    .B(\MuI._3155_ ),
    .Y(\MuI._3156_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4057_  (.A(\MuI._3037_ ),
    .B(\MuI._3156_ ),
    .Y(\MuI._3157_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4058_  (.A(\MuI._3082_ ),
    .B(\MuI._3083_ ),
    .X(\MuI._3158_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4059_  (.A1(\MuI._2994_ ),
    .A2(\MuI._3077_ ),
    .B1(\MuI._3078_ ),
    .Y(\MuI._3159_ ));
 sky130_fd_sc_hd__nand2_2 \MuI._4060_  (.A(\MuI._3079_ ),
    .B(\MuI._3159_ ),
    .Y(\MuI._3160_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4061_  (.A(\MuI._2905_ ),
    .B(\MuI._2879_ ),
    .C(\MuI._2904_ ),
    .X(\MuI._3161_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4062_  (.A(\MuI._0350_ ),
    .B(\MuI._2967_ ),
    .Y(\MuI._3162_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4063_  (.A1(\MuI._2887_ ),
    .A2(\MuI._3162_ ),
    .B1(\MuI._2968_ ),
    .X(\MuI._3163_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4064_  (.A1(\MuI._2905_ ),
    .A2(\MuI._2904_ ),
    .B1(\MuI._2879_ ),
    .Y(\MuI._3164_ ));
 sky130_fd_sc_hd__or3_2 \MuI._4065_  (.A(\MuI._3161_ ),
    .B(\MuI._3163_ ),
    .C(\MuI._3164_ ),
    .X(\MuI._3165_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4066_  (.A1(\MuI._3073_ ),
    .A2(\MuI._3074_ ),
    .B1(\MuI._3072_ ),
    .Y(\MuI._3166_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4067_  (.A(\MuI._3075_ ),
    .B(\MuI._3166_ ),
    .X(\MuI._3167_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4068_  (.A(\MuI._3165_ ),
    .B(\MuI._3167_ ),
    .X(\MuI._3168_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4069_  (.A(\MuI._2865_ ),
    .B(\MuI._2924_ ),
    .X(\MuI._3169_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4070_  (.A(\MuI._3165_ ),
    .B(\MuI._3167_ ),
    .Y(\MuI._3170_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4071_  (.A1(\MuI._3168_ ),
    .A2(\MuI._3169_ ),
    .B1(\MuI._3170_ ),
    .Y(\MuI._3171_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4072_  (.A(\MuI._3160_ ),
    .B(\MuI._3171_ ),
    .Y(\MuI._3172_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4073_  (.A(\MuI._2835_ ),
    .B(\MuI._2953_ ),
    .X(\MuI._3173_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4074_  (.A(\MuI._3160_ ),
    .B(\MuI._3171_ ),
    .Y(\MuI._3174_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4075_  (.A1(\MuI._3172_ ),
    .A2(\MuI._3173_ ),
    .B1(\MuI._3174_ ),
    .Y(\MuI._3175_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4076_  (.A(\MuI._3158_ ),
    .B(\MuI._3175_ ),
    .X(\MuI._3176_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4077_  (.A(\MuI._2418_ ),
    .B(\MuI._2958_ ),
    .Y(\MuI._3177_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4078_  (.A_N(\MuI._3175_ ),
    .B(\MuI._3158_ ),
    .X(\MuI._3178_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4079_  (.A1(\MuI._3176_ ),
    .A2(\MuI._3177_ ),
    .B1_N(\MuI._3178_ ),
    .X(\MuI._3179_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4080_  (.A(\MuI._3157_ ),
    .B(\MuI._3179_ ),
    .Y(\MuI._3180_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4081_  (.A(\MuI._2960_ ),
    .B(\MuI._3180_ ),
    .X(\MuI._3181_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4082_  (.A1(\MuI._2858_ ),
    .A2(\MuI._2859_ ),
    .B1(\MuI._2863_ ),
    .X(\MuI._3182_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4083_  (.A1(\MuI._2870_ ),
    .A2(\MuI._2877_ ),
    .B1(\MuI._2872_ ),
    .Y(\MuI._3183_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4084_  (.A1(\MuI._0570_ ),
    .A2(\MuI._2886_ ),
    .B1(\MuI._2882_ ),
    .B2(\MuI._0328_ ),
    .X(\MuI._3184_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4085_  (.A(\MuI._2880_ ),
    .X(\MuI._3185_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4086_  (.A(\MuI.a_operand[22] ),
    .B(\MuI._2894_ ),
    .C(\MuI._2892_ ),
    .D(\MuI._3185_ ),
    .X(\MuI._3186_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4087_  (.A1(\MuI._0801_ ),
    .A2(\MuI._2967_ ),
    .A3(\MuI._3184_ ),
    .B1(\MuI._3186_ ),
    .X(\MuI._3187_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4088_  (.A1(\MuI._2878_ ),
    .A2(\MuI._3183_ ),
    .B1(\MuI._3187_ ),
    .X(\MuI._3188_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4089_  (.A(\MuI.b_operand[7] ),
    .X(\MuI._3189_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4090_  (.A(\MuI.b_operand[6] ),
    .X(\MuI._3190_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4091_  (.A(\MuI.a_operand[19] ),
    .B(\MuI._1461_ ),
    .C(\MuI._3189_ ),
    .D(\MuI._3190_ ),
    .X(\MuI._3191_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4092_  (.A1(\MuI._1472_ ),
    .A2(\MuI._2867_ ),
    .B1(\MuI._2869_ ),
    .B2(\MuI._1010_ ),
    .Y(\MuI._3192_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4093_  (.A(\MuI._3191_ ),
    .B(\MuI._3192_ ),
    .Y(\MuI._3193_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4094_  (.A1(\MuI._2077_ ),
    .A2(\MuI._2898_ ),
    .A3(\MuI._3193_ ),
    .B1(\MuI._3191_ ),
    .X(\MuI._3194_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4095_  (.A(\MuI._2878_ ),
    .B(\MuI._3187_ ),
    .C(\MuI._3183_ ),
    .Y(\MuI._3195_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4096_  (.A1(\MuI._3188_ ),
    .A2(\MuI._3194_ ),
    .B1_N(\MuI._3195_ ),
    .X(\MuI._3196_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4097_  (.A1(\MuI._2864_ ),
    .A2(\MuI._3182_ ),
    .B1(\MuI._3196_ ),
    .X(\MuI._3197_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4098_  (.A(\MuI._2671_ ),
    .B(\MuI._2841_ ),
    .Y(\MuI._3198_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4099_  (.A1(\MuI._2605_ ),
    .A2(\MuI._2844_ ),
    .B1(\MuI._2845_ ),
    .B2(\MuI._2840_ ),
    .Y(\MuI._3199_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4100_  (.A(\MuI._2840_ ),
    .B(\MuI._2605_ ),
    .C(\MuI._2836_ ),
    .D(\MuI._2854_ ),
    .X(\MuI._3200_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4101_  (.A1(\MuI._3198_ ),
    .A2(\MuI._3199_ ),
    .B1_N(\MuI._3200_ ),
    .X(\MuI._3201_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4102_  (.A(\MuI._2616_ ),
    .B(\MuI._2850_ ),
    .Y(\MuI._3202_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4103_  (.A_N(\MuI._2856_ ),
    .B(\MuI._2855_ ),
    .X(\MuI._3203_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4104_  (.A(\MuI._3202_ ),
    .B(\MuI._3203_ ),
    .Y(\MuI._3204_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4105_  (.A_N(\MuI._3201_ ),
    .B(\MuI._3204_ ),
    .X(\MuI._3205_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4106_  (.A(\MuI._3204_ ),
    .B(\MuI._3201_ ),
    .Y(\MuI._3206_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4107_  (.A(\MuI._2804_ ),
    .B(\MuI._2801_ ),
    .Y(\MuI._3207_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4108_  (.A(\MuI._2798_ ),
    .B(\MuI._3207_ ),
    .Y(\MuI._3208_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4109_  (.A(\MuI._3206_ ),
    .B(\MuI._3208_ ),
    .X(\MuI._3209_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4110_  (.A(\MuI._3205_ ),
    .B(\MuI._3209_ ),
    .X(\MuI._3210_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4111_  (.A(\MuI._2864_ ),
    .B(\MuI._3196_ ),
    .C(\MuI._3182_ ),
    .Y(\MuI._3211_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4112_  (.A1(\MuI._3197_ ),
    .A2(\MuI._3210_ ),
    .B1_N(\MuI._3211_ ),
    .X(\MuI._3212_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4113_  (.A1(\MuI._2809_ ),
    .A2(\MuI._2810_ ),
    .B1(\MuI._2833_ ),
    .Y(\MuI._3213_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4114_  (.A(\MuI._2834_ ),
    .B(\MuI._3213_ ),
    .Y(\MuI._3214_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4115_  (.A(\MuI._3212_ ),
    .B(\MuI._3214_ ),
    .Y(\MuI._3215_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4116_  (.A(\MuI._2583_ ),
    .B(\MuI._2789_ ),
    .Y(\MuI._3216_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4117_  (.A1(\MuI._2919_ ),
    .A2(\MuI._2528_ ),
    .B1(\MuI._2539_ ),
    .B2(\MuI._2800_ ),
    .Y(\MuI._3217_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4118_  (.A(\MuI._2704_ ),
    .B(\MuI._2803_ ),
    .C(\MuI._2528_ ),
    .D(\MuI._2539_ ),
    .X(\MuI._3218_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4119_  (.A1(\MuI._3216_ ),
    .A2(\MuI._3217_ ),
    .B1_N(\MuI._3218_ ),
    .X(\MuI._3219_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4120_  (.A(\MuI._1274_ ),
    .B(\MuI._2787_ ),
    .Y(\MuI._3220_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4121_  (.A(\MuI._3220_ ),
    .B(\MuI._2793_ ),
    .Y(\MuI._3221_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4122_  (.A(\MuI._3219_ ),
    .B_N(\MuI._3221_ ),
    .X(\MuI._3222_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4123_  (.A(\MuI.a_operand[9] ),
    .X(\MuI._3223_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4124_  (.A(\MuI._3000_ ),
    .B(\MuI._2754_ ),
    .C(\MuI._2790_ ),
    .D(\MuI._3223_ ),
    .X(\MuI._3224_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4125_  (.A1(\MuI._1802_ ),
    .A2(\MuI._2773_ ),
    .B1(\MuI._2786_ ),
    .B2(\MuI._2550_ ),
    .Y(\MuI._3225_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4126_  (.A(\MuI._3224_ ),
    .B(\MuI._3225_ ),
    .Y(\MuI._3226_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4127_  (.A1(\MuI._1285_ ),
    .A2(\MuI._2363_ ),
    .A3(\MuI._3226_ ),
    .B1(\MuI._3224_ ),
    .X(\MuI._3227_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4128_  (.A(\MuI._3219_ ),
    .B(\MuI._3221_ ),
    .Y(\MuI._3228_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4129_  (.A(\MuI._3227_ ),
    .B(\MuI._3228_ ),
    .Y(\MuI._3229_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4130_  (.A(\MuI._2807_ ),
    .B(\MuI._2794_ ),
    .C(\MuI._2806_ ),
    .X(\MuI._3230_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4131_  (.A1(\MuI._2807_ ),
    .A2(\MuI._2806_ ),
    .B1(\MuI._2794_ ),
    .Y(\MuI._3231_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4132_  (.A(\MuI._3230_ ),
    .B(\MuI._3231_ ),
    .X(\MuI._3232_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4133_  (.A1(\MuI._3222_ ),
    .A2(\MuI._3229_ ),
    .B1(\MuI._3232_ ),
    .Y(\MuI._3233_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4134_  (.A(\MuI._3232_ ),
    .B(\MuI._3222_ ),
    .C(\MuI._3229_ ),
    .X(\MuI._3234_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4135_  (.A1_N(\MuI._0878_ ),
    .A2_N(\MuI._2385_ ),
    .B1(\MuI._2820_ ),
    .B2(\MuI._2821_ ),
    .X(\MuI._3235_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4136_  (.A(\MuI._2822_ ),
    .B(\MuI._3235_ ),
    .Y(\MuI._3236_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4137_  (.A(\MuI._0735_ ),
    .B(\MuI._2813_ ),
    .C(\MuI._2352_ ),
    .D(\MuI._2374_ ),
    .X(\MuI._3237_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4138_  (.A1(\MuI._1153_ ),
    .A2(\MuI._2363_ ),
    .B1(\MuI._2385_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._3238_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4139_  (.A_N(\MuI._3237_ ),
    .B_N(\MuI._3238_ ),
    .C(\MuI._2817_ ),
    .D(\MuI._2330_ ),
    .X(\MuI._3239_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4140_  (.A(\MuI._3237_ ),
    .B(\MuI._3239_ ),
    .Y(\MuI._3240_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4141_  (.A(\MuI._3236_ ),
    .B(\MuI._3240_ ),
    .Y(\MuI._3241_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4142_  (.A1(\MuI._0614_ ),
    .A2(\MuI._2330_ ),
    .B1(\MuI._2830_ ),
    .B2(\MuI._0361_ ),
    .Y(\MuI._3242_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4143_  (.A(\MuI._0361_ ),
    .B(\MuI._0614_ ),
    .C(\MuI._2330_ ),
    .D(\MuI._2830_ ),
    .X(\MuI._3243_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4144_  (.A(\MuI._3242_ ),
    .B(\MuI._3243_ ),
    .Y(\MuI._3244_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4145_  (.A(\MuI.a_operand[4] ),
    .X(\MuI._3245_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4146_  (.A(\MuI._3245_ ),
    .X(\MuI._3246_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4147_  (.A(\MuI._3246_ ),
    .X(\MuI._3247_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4148_  (.A(\MuI._3247_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._3248_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4149_  (.A(\MuI._3244_ ),
    .B(\MuI._3248_ ),
    .Y(\MuI._3249_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4150_  (.A(\MuI._3241_ ),
    .B(\MuI._3249_ ),
    .Y(\MuI._3250_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4151_  (.A(\MuI._3241_ ),
    .B(\MuI._3249_ ),
    .X(\MuI._3251_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4152_  (.A(\MuI._3250_ ),
    .B(\MuI._3251_ ),
    .Y(\MuI._3252_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4153_  (.A(\MuI._3233_ ),
    .B(\MuI._3234_ ),
    .C(\MuI._3252_ ),
    .Y(\MuI._3253_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4154_  (.A(\MuI._3233_ ),
    .B(\MuI._3253_ ),
    .X(\MuI._3254_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4155_  (.A(\MuI._3215_ ),
    .B(\MuI._3254_ ),
    .X(\MuI._3255_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4156_  (.A(\MuI._3211_ ),
    .B(\MuI._3197_ ),
    .Y(\MuI._3256_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4157_  (.A(\MuI._3256_ ),
    .B(\MuI._3210_ ),
    .Y(\MuI._3257_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4158_  (.A1(\MuI._3161_ ),
    .A2(\MuI._3164_ ),
    .B1(\MuI._3163_ ),
    .Y(\MuI._3258_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4159_  (.A(\MuI._3195_ ),
    .B(\MuI._3188_ ),
    .C(\MuI._3194_ ),
    .X(\MuI._3259_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4160_  (.A1(\MuI._3195_ ),
    .A2(\MuI._3188_ ),
    .B1(\MuI._3194_ ),
    .Y(\MuI._3260_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4161_  (.A(\MuI._3259_ ),
    .B(\MuI._3260_ ),
    .Y(\MuI._3261_ ));
 sky130_fd_sc_hd__buf_4 \MuI._4162_  (.A(\MuI.b_operand[1] ),
    .X(\MuI._3262_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4163_  (.A(\MuI.a_operand[22] ),
    .B(\MuI._3262_ ),
    .X(\MuI._3263_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4164_  (.A(\MuI._0570_ ),
    .B(\MuI._2886_ ),
    .Y(\MuI._3264_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4165_  (.A1(\MuI._3264_ ),
    .A2(\MuI._2883_ ),
    .B1(\MuI._3186_ ),
    .X(\MuI._3265_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4166_  (.A(\MuI._0790_ ),
    .B(\MuI._2967_ ),
    .Y(\MuI._3266_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4167_  (.A(\MuI._3265_ ),
    .B(\MuI._3266_ ),
    .X(\MuI._3267_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4168_  (.A(\MuI.b_operand[2] ),
    .X(\MuI._3268_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4169_  (.A(\MuI._3268_ ),
    .X(\MuI._3269_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._4170_  (.A1(\MuI._3263_ ),
    .A2(\MuI._3267_ ),
    .B1(\MuI._3269_ ),
    .C1(\MuI._0515_ ),
    .X(\MuI._3270_ ));
 sky130_fd_sc_hd__o22a_1 \MuI._4171_  (.A1(\MuI._2883_ ),
    .A2(\MuI._2887_ ),
    .B1(\MuI._2891_ ),
    .B2(\MuI._2893_ ),
    .X(\MuI._3271_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4172_  (.A(\MuI._2896_ ),
    .B(\MuI._3271_ ),
    .X(\MuI._3272_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4173_  (.A(\MuI._3270_ ),
    .B(\MuI._3272_ ),
    .X(\MuI._3273_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4174_  (.A(\MuI._3270_ ),
    .B(\MuI._3272_ ),
    .X(\MuI._3274_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4175_  (.A1(\MuI._3261_ ),
    .A2(\MuI._3273_ ),
    .B1(\MuI._3274_ ),
    .X(\MuI._3275_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4176_  (.A1(\MuI._3165_ ),
    .A2(\MuI._3258_ ),
    .B1(\MuI._3275_ ),
    .X(\MuI._3276_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4177_  (.A(\MuI._3165_ ),
    .B(\MuI._3275_ ),
    .C(\MuI._3258_ ),
    .X(\MuI._3277_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4178_  (.A1(\MuI._3257_ ),
    .A2(\MuI._3276_ ),
    .B1(\MuI._3277_ ),
    .Y(\MuI._3278_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4179_  (.A(\MuI._3168_ ),
    .B(\MuI._3169_ ),
    .Y(\MuI._3279_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4180_  (.A(\MuI._3278_ ),
    .B(\MuI._3279_ ),
    .X(\MuI._3280_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4181_  (.A(\MuI._3278_ ),
    .B(\MuI._3279_ ),
    .Y(\MuI._3281_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4182_  (.A1(\MuI._3255_ ),
    .A2(\MuI._3280_ ),
    .B1(\MuI._3281_ ),
    .Y(\MuI._3282_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4183_  (.A(\MuI._3160_ ),
    .B(\MuI._3171_ ),
    .Y(\MuI._3283_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4184_  (.A(\MuI._3283_ ),
    .B(\MuI._3173_ ),
    .Y(\MuI._3284_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4185_  (.A_N(\MuI._3282_ ),
    .B(\MuI._3284_ ),
    .X(\MuI._3285_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4186_  (.A(\MuI._2834_ ),
    .B(\MuI._3212_ ),
    .C(\MuI._3213_ ),
    .X(\MuI._3286_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4187_  (.A1(\MuI._3215_ ),
    .A2(\MuI._3254_ ),
    .B1(\MuI._3286_ ),
    .Y(\MuI._3287_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4188_  (.A(\MuI._2824_ ),
    .B(\MuI._2832_ ),
    .Y(\MuI._3288_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._4189_  (.A1(\MuI._2816_ ),
    .A2(\MuI._2818_ ),
    .A3(\MuI._2823_ ),
    .B1(\MuI._3288_ ),
    .X(\MuI._3289_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4190_  (.A(\MuI._3287_ ),
    .B(\MuI._3289_ ),
    .X(\MuI._3290_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4191_  (.A1(\MuI._2825_ ),
    .A2(\MuI._2831_ ),
    .B1_N(\MuI._2827_ ),
    .X(\MuI._3291_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4192_  (.A(\MuI._3290_ ),
    .B(\MuI._3291_ ),
    .Y(\MuI._3292_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4193_  (.A(\MuI._3282_ ),
    .B(\MuI._3284_ ),
    .Y(\MuI._3293_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4194_  (.A(\MuI._3292_ ),
    .B(\MuI._3293_ ),
    .X(\MuI._3294_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4195_  (.A(\MuI._3176_ ),
    .B(\MuI._3177_ ),
    .X(\MuI._3295_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4196_  (.A1(\MuI._3285_ ),
    .A2(\MuI._3294_ ),
    .B1(\MuI._3295_ ),
    .Y(\MuI._3296_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4197_  (.A(\MuI._3285_ ),
    .B(\MuI._3294_ ),
    .C(\MuI._3295_ ),
    .X(\MuI._3297_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4198_  (.A(\MuI._3296_ ),
    .B(\MuI._3297_ ),
    .Y(\MuI._3298_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4199_  (.A(\MuI._3291_ ),
    .B_N(\MuI._3290_ ),
    .X(\MuI._3299_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._4200_  (.A1(\MuI._3287_ ),
    .A2(\MuI._3289_ ),
    .B1(\MuI._3299_ ),
    .Y(\MuI._3300_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4201_  (.A(\MuI._3298_ ),
    .B_N(\MuI._3300_ ),
    .X(\MuI._3301_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4202_  (.A(\MuI._3181_ ),
    .B(\MuI._3296_ ),
    .C(\MuI._3301_ ),
    .X(\MuI._3302_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4203_  (.A1(\MuI._3296_ ),
    .A2(\MuI._3301_ ),
    .B1(\MuI._3181_ ),
    .X(\MuI._3303_ ));
 sky130_fd_sc_hd__nor2b_1 \MuI._4204_  (.A(\MuI._3302_ ),
    .B_N(\MuI._3303_ ),
    .Y(\MuI._3304_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4205_  (.A(\MuI._3300_ ),
    .B(\MuI._3298_ ),
    .X(\MuI._3305_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4206_  (.A(\MuI.b_operand[4] ),
    .X(\MuI._3306_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4207_  (.A(\MuI.b_operand[3] ),
    .X(\MuI._3307_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4208_  (.A(\MuI._0559_ ),
    .B(\MuI.a_operand[20] ),
    .C(\MuI._3306_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._3308_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4209_  (.A1(\MuI._0768_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._3185_ ),
    .B2(\MuI._0559_ ),
    .Y(\MuI._3309_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4210_  (.A(\MuI._3308_ ),
    .B(\MuI._3309_ ),
    .X(\MuI._3310_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4211_  (.A(\MuI._1021_ ),
    .B(\MuI._2895_ ),
    .Y(\MuI._3311_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4212_  (.A(\MuI._3310_ ),
    .B(\MuI._3311_ ),
    .Y(\MuI._3312_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4213_  (.A(\MuI._2843_ ),
    .B(\MuI._2871_ ),
    .Y(\MuI._3313_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4214_  (.A(\MuI._3313_ ),
    .B(\MuI._3193_ ),
    .Y(\MuI._3314_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4215_  (.A1(\MuI._3308_ ),
    .A2(\MuI._3312_ ),
    .B1(\MuI._3314_ ),
    .Y(\MuI._3315_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4216_  (.A(\MuI._3091_ ),
    .B(\MuI._2898_ ),
    .Y(\MuI._3316_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4217_  (.A1(\MuI._2066_ ),
    .A2(\MuI._2874_ ),
    .B1(\MuI._2876_ ),
    .B2(\MuI._1483_ ),
    .Y(\MuI._3317_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4218_  (.A(\MuI._1472_ ),
    .B(\MuI._2843_ ),
    .C(\MuI._2874_ ),
    .D(\MuI._2876_ ),
    .X(\MuI._3318_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4219_  (.A1(\MuI._3316_ ),
    .A2(\MuI._3317_ ),
    .B1_N(\MuI._3318_ ),
    .X(\MuI._3319_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4220_  (.A(\MuI._3308_ ),
    .B(\MuI._3312_ ),
    .C(\MuI._3314_ ),
    .X(\MuI._3320_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4221_  (.A(\MuI._3315_ ),
    .B(\MuI._3320_ ),
    .X(\MuI._3321_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4222_  (.A(\MuI._3319_ ),
    .B_N(\MuI._3321_ ),
    .X(\MuI._3322_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4223_  (.A(\MuI._3206_ ),
    .B(\MuI._3208_ ),
    .Y(\MuI._3323_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4224_  (.A(\MuI._3209_ ),
    .B(\MuI._3323_ ),
    .X(\MuI._3324_ ));
 sky130_fd_sc_hd__a21o_2 \MuI._4225_  (.A1(\MuI._3315_ ),
    .A2(\MuI._3322_ ),
    .B1(\MuI._3324_ ),
    .X(\MuI._3325_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4226_  (.A(\MuI._2528_ ),
    .B(\MuI._2850_ ),
    .Y(\MuI._3326_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4227_  (.A1(\MuI._2671_ ),
    .A2(\MuI._2975_ ),
    .B1(\MuI._2976_ ),
    .B2(\MuI._2616_ ),
    .Y(\MuI._3327_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4228_  (.A(\MuI._2616_ ),
    .B(\MuI._2660_ ),
    .C(\MuI._2844_ ),
    .D(\MuI._2845_ ),
    .X(\MuI._3328_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4229_  (.A1(\MuI._3326_ ),
    .A2(\MuI._3327_ ),
    .B1_N(\MuI._3328_ ),
    .X(\MuI._3329_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4230_  (.A(\MuI._3200_ ),
    .B(\MuI._3199_ ),
    .Y(\MuI._3330_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4231_  (.A(\MuI._3198_ ),
    .B(\MuI._3330_ ),
    .Y(\MuI._3331_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4232_  (.A_N(\MuI._3329_ ),
    .B(\MuI._3331_ ),
    .X(\MuI._3332_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4233_  (.A(\MuI._3331_ ),
    .B(\MuI._3329_ ),
    .Y(\MuI._3333_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4234_  (.A(\MuI._3218_ ),
    .B(\MuI._3217_ ),
    .Y(\MuI._3334_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4235_  (.A(\MuI._3216_ ),
    .B(\MuI._3334_ ),
    .Y(\MuI._3335_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4236_  (.A(\MuI._3333_ ),
    .B(\MuI._3335_ ),
    .X(\MuI._3336_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4237_  (.A(\MuI._3315_ ),
    .B(\MuI._3322_ ),
    .C(\MuI._3324_ ),
    .Y(\MuI._3337_ ));
 sky130_fd_sc_hd__o211ai_4 \MuI._4238_  (.A1(\MuI._3332_ ),
    .A2(\MuI._3336_ ),
    .B1(\MuI._3325_ ),
    .C1(\MuI._3337_ ),
    .Y(\MuI._3338_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4239_  (.A1(\MuI._3233_ ),
    .A2(\MuI._3234_ ),
    .B1(\MuI._3252_ ),
    .X(\MuI._3339_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._4240_  (.A1(\MuI._3325_ ),
    .A2(\MuI._3338_ ),
    .B1(\MuI._3339_ ),
    .C1(\MuI._3253_ ),
    .Y(\MuI._3340_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4241_  (.A1(\MuI._3253_ ),
    .A2(\MuI._3339_ ),
    .B1(\MuI._3338_ ),
    .C1(\MuI._3325_ ),
    .Y(\MuI._3341_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4242_  (.A(\MuI._2796_ ),
    .B(\MuI._2791_ ),
    .Y(\MuI._3342_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4243_  (.A1(\MuI._2919_ ),
    .A2(\MuI._2539_ ),
    .B1(\MuI._2789_ ),
    .B2(\MuI._2800_ ),
    .Y(\MuI._3343_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4244_  (.A(\MuI._2704_ ),
    .B(\MuI._2803_ ),
    .C(\MuI._2539_ ),
    .D(\MuI._2495_ ),
    .X(\MuI._3344_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4245_  (.A1(\MuI._3342_ ),
    .A2(\MuI._3343_ ),
    .B1_N(\MuI._3344_ ),
    .X(\MuI._3345_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4246_  (.A(\MuI._2473_ ),
    .B(\MuI._2363_ ),
    .Y(\MuI._3346_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4247_  (.A(\MuI._3346_ ),
    .B(\MuI._3226_ ),
    .Y(\MuI._3347_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4248_  (.A(\MuI._3345_ ),
    .B_N(\MuI._3347_ ),
    .X(\MuI._3348_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4249_  (.A(\MuI.a_operand[8] ),
    .X(\MuI._3349_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4250_  (.A(\MuI._3000_ ),
    .B(\MuI._2754_ ),
    .C(\MuI._3223_ ),
    .D(\MuI._3349_ ),
    .X(\MuI._3350_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4251_  (.A1(\MuI._2517_ ),
    .A2(\MuI._2786_ ),
    .B1(\MuI._2352_ ),
    .B2(\MuI._2550_ ),
    .Y(\MuI._3351_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4252_  (.A(\MuI._3350_ ),
    .B(\MuI._3351_ ),
    .Y(\MuI._3352_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4253_  (.A1(\MuI._1285_ ),
    .A2(\MuI._2385_ ),
    .A3(\MuI._3352_ ),
    .B1(\MuI._3350_ ),
    .X(\MuI._3353_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4254_  (.A(\MuI._3345_ ),
    .B(\MuI._3347_ ),
    .Y(\MuI._3354_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4255_  (.A(\MuI._3353_ ),
    .B(\MuI._3354_ ),
    .Y(\MuI._3355_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4256_  (.A(\MuI._3227_ ),
    .B(\MuI._3228_ ),
    .Y(\MuI._3356_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4257_  (.A1(\MuI._3348_ ),
    .A2(\MuI._3355_ ),
    .B1(\MuI._3356_ ),
    .Y(\MuI._3357_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4258_  (.A(\MuI._3348_ ),
    .B(\MuI._3355_ ),
    .C(\MuI._3356_ ),
    .X(\MuI._3358_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4259_  (.A1_N(\MuI._2817_ ),
    .A2_N(\MuI._2330_ ),
    .B1(\MuI._3237_ ),
    .B2(\MuI._3238_ ),
    .X(\MuI._3359_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4260_  (.A(\MuI._3239_ ),
    .B(\MuI._3359_ ),
    .Y(\MuI._3360_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4261_  (.A(\MuI.b_operand[20] ),
    .B(\MuI._2830_ ),
    .Y(\MuI._3361_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4262_  (.A(\MuI.a_operand[6] ),
    .X(\MuI._3362_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4263_  (.A(\MuI._3362_ ),
    .X(\MuI._3363_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4264_  (.A1(\MuI._1142_ ),
    .A2(\MuI._2374_ ),
    .B1(\MuI._3363_ ),
    .B2(\MuI._2939_ ),
    .Y(\MuI._3364_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4265_  (.A(\MuI.b_operand[19] ),
    .B(\MuI._2811_ ),
    .C(\MuI._2374_ ),
    .D(\MuI._2319_ ),
    .X(\MuI._3365_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4266_  (.A1(\MuI._3361_ ),
    .A2(\MuI._3364_ ),
    .B1_N(\MuI._3365_ ),
    .X(\MuI._3366_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4267_  (.A(\MuI._3360_ ),
    .B(\MuI._3366_ ),
    .Y(\MuI._3367_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4268_  (.A1(\MuI._0614_ ),
    .A2(\MuI._2830_ ),
    .B1(\MuI._3247_ ),
    .B2(\MuI._0361_ ),
    .Y(\MuI._3368_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4269_  (.A(\MuI._0361_ ),
    .B(\MuI._0614_ ),
    .C(\MuI._2830_ ),
    .D(\MuI._3247_ ),
    .X(\MuI._3369_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4270_  (.A(\MuI._3368_ ),
    .B(\MuI._3369_ ),
    .Y(\MuI._3370_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4271_  (.A(\MuI.a_operand[3] ),
    .X(\MuI._3371_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4272_  (.A(\MuI._3371_ ),
    .X(\MuI._3372_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4273_  (.A(\MuI._3372_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._3373_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4274_  (.A(\MuI._3370_ ),
    .B(\MuI._3373_ ),
    .Y(\MuI._3374_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4275_  (.A(\MuI._3367_ ),
    .B(\MuI._3374_ ),
    .Y(\MuI._3375_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4276_  (.A(\MuI._3367_ ),
    .B(\MuI._3374_ ),
    .X(\MuI._3376_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4277_  (.A(\MuI._3375_ ),
    .B(\MuI._3376_ ),
    .Y(\MuI._3377_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4278_  (.A(\MuI._3357_ ),
    .B(\MuI._3358_ ),
    .C(\MuI._3377_ ),
    .Y(\MuI._3378_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4279_  (.A(\MuI._3357_ ),
    .B(\MuI._3378_ ),
    .X(\MuI._3379_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._4280_  (.A_N(\MuI._3340_ ),
    .B(\MuI._3341_ ),
    .C(\MuI._3379_ ),
    .X(\MuI._3380_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._4281_  (.A1(\MuI._2822_ ),
    .A2(\MuI._3235_ ),
    .A3(\MuI._3240_ ),
    .B1(\MuI._3250_ ),
    .X(\MuI._3381_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._4282_  (.A1(\MuI._3340_ ),
    .A2(\MuI._3380_ ),
    .B1_N(\MuI._3381_ ),
    .Y(\MuI._3382_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4283_  (.A1(\MuI._3242_ ),
    .A2(\MuI._3248_ ),
    .B1_N(\MuI._3243_ ),
    .X(\MuI._3383_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._4284_  (.A(\MuI._3340_ ),
    .B(\MuI._3380_ ),
    .C_N(\MuI._3381_ ),
    .X(\MuI._3384_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4285_  (.A(\MuI._3382_ ),
    .B(\MuI._3384_ ),
    .X(\MuI._3385_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4286_  (.A(\MuI._3383_ ),
    .B_N(\MuI._3385_ ),
    .X(\MuI._3386_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4287_  (.A(\MuI._3382_ ),
    .B(\MuI._3386_ ),
    .Y(\MuI._3387_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4288_  (.A(\MuI._3385_ ),
    .B(\MuI._3383_ ),
    .Y(\MuI._3388_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4289_  (.A(\MuI._3340_ ),
    .B_N(\MuI._3341_ ),
    .X(\MuI._3389_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4290_  (.A(\MuI._3389_ ),
    .B(\MuI._3379_ ),
    .Y(\MuI._3390_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4291_  (.A1(\MuI._3325_ ),
    .A2(\MuI._3337_ ),
    .B1(\MuI._3332_ ),
    .C1(\MuI._3336_ ),
    .X(\MuI._3391_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4292_  (.A(\MuI._3338_ ),
    .B(\MuI._3391_ ),
    .X(\MuI._3392_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4293_  (.A(\MuI._3321_ ),
    .B(\MuI._3319_ ),
    .Y(\MuI._3393_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4294_  (.A(\MuI._3310_ ),
    .B(\MuI._3311_ ),
    .X(\MuI._3394_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4295_  (.A(\MuI._3312_ ),
    .B(\MuI._3394_ ),
    .Y(\MuI._3395_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4296_  (.A(\MuI.b_operand[0] ),
    .X(\MuI._3396_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4297_  (.A(\MuI._3396_ ),
    .X(\MuI._3397_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._4298_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._3397_ ),
    .X(\MuI._3398_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4299_  (.A(\MuI._3263_ ),
    .B(\MuI._3398_ ),
    .X(\MuI._3399_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4300_  (.A(\MuI._3263_ ),
    .B(\MuI._3398_ ),
    .X(\MuI._3400_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4301_  (.A1(\MuI._0570_ ),
    .A2(\MuI._3269_ ),
    .A3(\MuI._3399_ ),
    .B1(\MuI._3400_ ),
    .X(\MuI._3401_ ));
 sky130_fd_sc_hd__buf_4 \MuI._4302_  (.A(\MuI.b_operand[1] ),
    .X(\MuI._3402_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4303_  (.A(\MuI._3402_ ),
    .X(\MuI._3403_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4304_  (.A1(\MuI._0339_ ),
    .A2(\MuI._3269_ ),
    .B1(\MuI._3403_ ),
    .B2(\MuI._0504_ ),
    .Y(\MuI._3404_ ));
 sky130_fd_sc_hd__a31oi_2 \MuI._4305_  (.A1(\MuI._3269_ ),
    .A2(\MuI._0504_ ),
    .A3(\MuI._3263_ ),
    .B1(\MuI._3404_ ),
    .Y(\MuI._3405_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4306_  (.A(\MuI._3401_ ),
    .B(\MuI._3405_ ),
    .X(\MuI._3406_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4307_  (.A(\MuI._3401_ ),
    .B(\MuI._3405_ ),
    .Y(\MuI._3407_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4308_  (.A1(\MuI._3395_ ),
    .A2(\MuI._3406_ ),
    .B1_N(\MuI._3407_ ),
    .X(\MuI._3408_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._4309_  (.A_N(\MuI._3263_ ),
    .B(\MuI._3269_ ),
    .C(\MuI._0515_ ),
    .X(\MuI._3409_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4310_  (.A(\MuI._3267_ ),
    .B(\MuI._3409_ ),
    .Y(\MuI._3410_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4311_  (.A(\MuI._3408_ ),
    .B(\MuI._3410_ ),
    .Y(\MuI._3411_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4312_  (.A_N(\MuI._3410_ ),
    .B(\MuI._3408_ ),
    .X(\MuI._3412_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4313_  (.A1(\MuI._3393_ ),
    .A2(\MuI._3411_ ),
    .B1(\MuI._3412_ ),
    .X(\MuI._3413_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4314_  (.A(\MuI._3274_ ),
    .B_N(\MuI._3273_ ),
    .X(\MuI._3414_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4315_  (.A(\MuI._3261_ ),
    .B(\MuI._3414_ ),
    .Y(\MuI._3415_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4316_  (.A(\MuI._3413_ ),
    .B(\MuI._3415_ ),
    .X(\MuI._3416_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4317_  (.A(\MuI._3413_ ),
    .B(\MuI._3415_ ),
    .X(\MuI._3417_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4318_  (.A1(\MuI._3392_ ),
    .A2(\MuI._3416_ ),
    .B1(\MuI._3417_ ),
    .Y(\MuI._3418_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4319_  (.A_N(\MuI._3277_ ),
    .B(\MuI._3276_ ),
    .X(\MuI._3419_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4320_  (.A(\MuI._3257_ ),
    .B(\MuI._3419_ ),
    .X(\MuI._3420_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4321_  (.A(\MuI._3418_ ),
    .B(\MuI._3420_ ),
    .Y(\MuI._3421_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4322_  (.A_N(\MuI._3418_ ),
    .B(\MuI._3420_ ),
    .X(\MuI._3422_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4323_  (.A1(\MuI._3390_ ),
    .A2(\MuI._3421_ ),
    .B1(\MuI._3422_ ),
    .Y(\MuI._0000_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4324_  (.A(\MuI._3255_ ),
    .B(\MuI._3280_ ),
    .X(\MuI._0001_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4325_  (.A(\MuI._3255_ ),
    .B(\MuI._3280_ ),
    .Y(\MuI._0002_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4326_  (.A(\MuI._0001_ ),
    .B(\MuI._0002_ ),
    .Y(\MuI._0003_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4327_  (.A(\MuI._0000_ ),
    .B(\MuI._0003_ ),
    .Y(\MuI._0004_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4328_  (.A(\MuI._0001_ ),
    .B(\MuI._0000_ ),
    .C(\MuI._0002_ ),
    .X(\MuI._0005_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4329_  (.A1(\MuI._3388_ ),
    .A2(\MuI._0004_ ),
    .B1_N(\MuI._0005_ ),
    .Y(\MuI._0006_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4330_  (.A(\MuI._3292_ ),
    .B(\MuI._3293_ ),
    .Y(\MuI._0007_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4331_  (.A(\MuI._3294_ ),
    .B(\MuI._0007_ ),
    .X(\MuI._0008_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4332_  (.A(\MuI._0006_ ),
    .B(\MuI._0008_ ),
    .X(\MuI._0009_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4333_  (.A(\MuI._0006_ ),
    .B(\MuI._0008_ ),
    .Y(\MuI._0011_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4334_  (.A1(\MuI._3387_ ),
    .A2(\MuI._0009_ ),
    .B1(\MuI._0011_ ),
    .Y(\MuI._0012_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4335_  (.A(\MuI._3305_ ),
    .B(\MuI._0012_ ),
    .X(\MuI._0013_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4336_  (.A(\MuI._3304_ ),
    .B(\MuI._0013_ ),
    .Y(\MuI._0014_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4337_  (.A(\MuI._3387_ ),
    .B(\MuI._0009_ ),
    .Y(\MuI._0015_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4338_  (.A(\MuI._3388_ ),
    .B(\MuI._0004_ ),
    .Y(\MuI._0016_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4339_  (.A(\MuI.b_operand[1] ),
    .X(\MuI._0017_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4340_  (.A(\MuI.b_operand[0] ),
    .X(\MuI._0018_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4341_  (.A(\MuI.a_operand[22] ),
    .B(\MuI._0559_ ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._0019_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4342_  (.A(\MuI._0018_ ),
    .X(\MuI._0020_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4343_  (.A1(\MuI._0559_ ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI.a_operand[22] ),
    .Y(\MuI._0022_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4344_  (.A_N(\MuI._0019_ ),
    .B_N(\MuI._0022_ ),
    .C(\MuI._0768_ ),
    .D(\MuI._3268_ ),
    .X(\MuI._0023_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4345_  (.A(\MuI._0019_ ),
    .B(\MuI._0023_ ),
    .X(\MuI._0024_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4346_  (.A(\MuI._0570_ ),
    .B(\MuI._3269_ ),
    .Y(\MuI._0025_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4347_  (.A(\MuI._0025_ ),
    .B(\MuI._3399_ ),
    .Y(\MuI._0026_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4348_  (.A(\MuI._0024_ ),
    .B(\MuI._0026_ ),
    .X(\MuI._0027_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4349_  (.A(\MuI._1494_ ),
    .B(\MuI._2967_ ),
    .Y(\MuI._0028_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4350_  (.A1(\MuI._1032_ ),
    .A2(\MuI._2886_ ),
    .B1(\MuI._2882_ ),
    .B2(\MuI._0790_ ),
    .Y(\MuI._0029_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4351_  (.A(\MuI._0790_ ),
    .B(\MuI._1021_ ),
    .C(\MuI._2886_ ),
    .D(\MuI._2882_ ),
    .X(\MuI._0030_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4352_  (.A(\MuI._0029_ ),
    .B(\MuI._0030_ ),
    .Y(\MuI._0031_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4353_  (.A(\MuI._0028_ ),
    .B(\MuI._0031_ ),
    .Y(\MuI._0033_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4354_  (.A(\MuI._0024_ ),
    .B(\MuI._0026_ ),
    .X(\MuI._0034_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4355_  (.A1(\MuI._0027_ ),
    .A2(\MuI._0033_ ),
    .B1(\MuI._0034_ ),
    .Y(\MuI._0035_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4356_  (.A(\MuI._3395_ ),
    .B(\MuI._3406_ ),
    .Y(\MuI._0036_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4357_  (.A(\MuI._0035_ ),
    .B(\MuI._0036_ ),
    .X(\MuI._0037_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4358_  (.A(\MuI._2616_ ),
    .B(\MuI._2871_ ),
    .Y(\MuI._0038_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4359_  (.A1(\MuI._2840_ ),
    .A2(\MuI._2867_ ),
    .B1(\MuI._2869_ ),
    .B2(\MuI._2843_ ),
    .Y(\MuI._0039_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4360_  (.A(\MuI._2055_ ),
    .B(\MuI._2852_ ),
    .C(\MuI._2873_ ),
    .D(\MuI._2875_ ),
    .X(\MuI._0040_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4361_  (.A1(\MuI._0038_ ),
    .A2(\MuI._0039_ ),
    .B1_N(\MuI._0040_ ),
    .X(\MuI._0041_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4362_  (.A1(\MuI._0028_ ),
    .A2(\MuI._0029_ ),
    .B1_N(\MuI._0030_ ),
    .X(\MuI._0042_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4363_  (.A(\MuI._3318_ ),
    .B(\MuI._3317_ ),
    .Y(\MuI._0044_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4364_  (.A(\MuI._3316_ ),
    .B(\MuI._0044_ ),
    .Y(\MuI._0045_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4365_  (.A(\MuI._0042_ ),
    .B(\MuI._0045_ ),
    .Y(\MuI._0046_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4366_  (.A(\MuI._0041_ ),
    .B(\MuI._0046_ ),
    .Y(\MuI._0047_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4367_  (.A(\MuI._0035_ ),
    .B(\MuI._0036_ ),
    .Y(\MuI._0048_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4368_  (.A1(\MuI._0037_ ),
    .A2(\MuI._0047_ ),
    .B1(\MuI._0048_ ),
    .Y(\MuI._0049_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4369_  (.A(\MuI._3393_ ),
    .B(\MuI._3411_ ),
    .X(\MuI._0050_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4370_  (.A(\MuI._0049_ ),
    .B(\MuI._0050_ ),
    .Y(\MuI._0051_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4371_  (.A(\MuI._2850_ ),
    .B(\MuI._2539_ ),
    .Y(\MuI._0052_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4372_  (.A1(\MuI._2440_ ),
    .A2(\MuI._2975_ ),
    .B1(\MuI._2976_ ),
    .B2(\MuI._2671_ ),
    .Y(\MuI._0053_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4373_  (.A(\MuI._2660_ ),
    .B(\MuI._2440_ ),
    .C(\MuI._2844_ ),
    .D(\MuI._2845_ ),
    .X(\MuI._0055_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4374_  (.A1(\MuI._0052_ ),
    .A2(\MuI._0053_ ),
    .B1_N(\MuI._0055_ ),
    .X(\MuI._0056_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4375_  (.A(\MuI._3328_ ),
    .B(\MuI._3327_ ),
    .Y(\MuI._0057_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4376_  (.A(\MuI._3326_ ),
    .B(\MuI._0057_ ),
    .Y(\MuI._0058_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4377_  (.A(\MuI._0056_ ),
    .B_N(\MuI._0058_ ),
    .X(\MuI._0059_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4378_  (.A(\MuI._0058_ ),
    .B(\MuI._0056_ ),
    .Y(\MuI._0060_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4379_  (.A(\MuI._3344_ ),
    .B(\MuI._3343_ ),
    .Y(\MuI._0061_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4380_  (.A(\MuI._3342_ ),
    .B(\MuI._0061_ ),
    .Y(\MuI._0062_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4381_  (.A(\MuI._0060_ ),
    .B(\MuI._0062_ ),
    .Y(\MuI._0063_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4382_  (.A(\MuI._0042_ ),
    .B_N(\MuI._0045_ ),
    .X(\MuI._0064_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4383_  (.A(\MuI._0041_ ),
    .B_N(\MuI._0046_ ),
    .X(\MuI._0066_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4384_  (.A(\MuI._3333_ ),
    .B(\MuI._3335_ ),
    .Y(\MuI._0067_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4385_  (.A(\MuI._3336_ ),
    .B(\MuI._0067_ ),
    .X(\MuI._0068_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4386_  (.A1(\MuI._0064_ ),
    .A2(\MuI._0066_ ),
    .B1(\MuI._0068_ ),
    .Y(\MuI._0069_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4387_  (.A(\MuI._0064_ ),
    .B(\MuI._0066_ ),
    .C(\MuI._0068_ ),
    .X(\MuI._0070_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4388_  (.A1(\MuI._0059_ ),
    .A2(\MuI._0063_ ),
    .B1(\MuI._0069_ ),
    .C1(\MuI._0070_ ),
    .X(\MuI._0071_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4389_  (.A1(\MuI._0069_ ),
    .A2(\MuI._0070_ ),
    .B1(\MuI._0059_ ),
    .C1(\MuI._0063_ ),
    .Y(\MuI._0072_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4390_  (.A(\MuI._0071_ ),
    .B(\MuI._0072_ ),
    .X(\MuI._0073_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4391_  (.A_N(\MuI._0049_ ),
    .B(\MuI._0050_ ),
    .X(\MuI._0074_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._4392_  (.A1(\MuI._0051_ ),
    .A2(\MuI._0073_ ),
    .B1(\MuI._0074_ ),
    .Y(\MuI._0075_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4393_  (.A(\MuI._3392_ ),
    .B(\MuI._3416_ ),
    .Y(\MuI._0076_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4394_  (.A(\MuI._0075_ ),
    .B(\MuI._0076_ ),
    .X(\MuI._0077_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4395_  (.A(\MuI._2796_ ),
    .B(\MuI._2786_ ),
    .Y(\MuI._0078_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4396_  (.A1(\MuI._2919_ ),
    .A2(\MuI._2495_ ),
    .B1(\MuI._2791_ ),
    .B2(\MuI._2800_ ),
    .Y(\MuI._0079_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4397_  (.A(\MuI._2704_ ),
    .B(\MuI._2649_ ),
    .C(\MuI._2495_ ),
    .D(\MuI._2773_ ),
    .X(\MuI._0080_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4398_  (.A1(\MuI._0078_ ),
    .A2(\MuI._0079_ ),
    .B1_N(\MuI._0080_ ),
    .X(\MuI._0081_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4399_  (.A(\MuI._2473_ ),
    .B(\MuI._2374_ ),
    .Y(\MuI._0082_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4400_  (.A(\MuI._0082_ ),
    .B(\MuI._3352_ ),
    .Y(\MuI._0083_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4401_  (.A(\MuI._0081_ ),
    .B_N(\MuI._0083_ ),
    .X(\MuI._0084_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4402_  (.A(\MuI.a_operand[7] ),
    .X(\MuI._0085_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4403_  (.A(\MuI._1296_ ),
    .B(\MuI.b_operand[15] ),
    .C(\MuI._2341_ ),
    .D(\MuI._0085_ ),
    .X(\MuI._0087_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4404_  (.A(\MuI.a_operand[7] ),
    .X(\MuI._0088_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4405_  (.A1(\MuI._1791_ ),
    .A2(\MuI._3349_ ),
    .B1(\MuI._0088_ ),
    .B2(\MuI._3000_ ),
    .Y(\MuI._0089_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4406_  (.A_N(\MuI._0087_ ),
    .B_N(\MuI._0089_ ),
    .C(\MuI.b_operand[17] ),
    .D(\MuI._3363_ ),
    .X(\MuI._0090_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4407_  (.A(\MuI._0081_ ),
    .B(\MuI._0083_ ),
    .Y(\MuI._0091_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4408_  (.A1(\MuI._0087_ ),
    .A2(\MuI._0090_ ),
    .B1(\MuI._0091_ ),
    .Y(\MuI._0092_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4409_  (.A(\MuI._3353_ ),
    .B(\MuI._3354_ ),
    .Y(\MuI._0093_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4410_  (.A1(\MuI._0084_ ),
    .A2(\MuI._0092_ ),
    .B1(\MuI._0093_ ),
    .Y(\MuI._0094_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4411_  (.A(\MuI._0084_ ),
    .B(\MuI._0092_ ),
    .C(\MuI._0093_ ),
    .X(\MuI._0095_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4412_  (.A(\MuI._3365_ ),
    .B(\MuI._3364_ ),
    .Y(\MuI._0096_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4413_  (.A(\MuI._3361_ ),
    .B(\MuI._0096_ ),
    .Y(\MuI._0098_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4414_  (.A(\MuI.b_operand[20] ),
    .B(\MuI._3247_ ),
    .Y(\MuI._0099_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4415_  (.A(\MuI.a_operand[5] ),
    .X(\MuI._0100_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4416_  (.A(\MuI._0100_ ),
    .X(\MuI._0101_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4417_  (.A1(\MuI._2813_ ),
    .A2(\MuI._3363_ ),
    .B1(\MuI._0101_ ),
    .B2(\MuI._2814_ ),
    .Y(\MuI._0102_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4418_  (.A(\MuI._2939_ ),
    .B(\MuI._2811_ ),
    .C(\MuI._3363_ ),
    .D(\MuI._0101_ ),
    .X(\MuI._0103_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4419_  (.A1(\MuI._0099_ ),
    .A2(\MuI._0102_ ),
    .B1_N(\MuI._0103_ ),
    .X(\MuI._0104_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4420_  (.A(\MuI._0098_ ),
    .B(\MuI._0104_ ),
    .Y(\MuI._0105_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4421_  (.A1(\MuI.b_operand[21] ),
    .A2(\MuI._3247_ ),
    .B1(\MuI._3372_ ),
    .B2(\MuI._2826_ ),
    .Y(\MuI._0106_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4422_  (.A(\MuI.b_operand[22] ),
    .B(\MuI.b_operand[21] ),
    .C(\MuI._3247_ ),
    .D(\MuI._3372_ ),
    .X(\MuI._0107_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4423_  (.A(\MuI._0106_ ),
    .B(\MuI._0107_ ),
    .Y(\MuI._0109_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4424_  (.A(\MuI.a_operand[2] ),
    .X(\MuI._0110_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4425_  (.A(\MuI._0110_ ),
    .X(\MuI._0111_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4426_  (.A(\MuI._0111_ ),
    .X(\MuI._0112_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4427_  (.A(\MuI._0112_ ),
    .B(\MuI._0438_ ),
    .Y(\MuI._0113_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4428_  (.A(\MuI._0109_ ),
    .B(\MuI._0113_ ),
    .Y(\MuI._0114_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4429_  (.A(\MuI._0105_ ),
    .B(\MuI._0114_ ),
    .X(\MuI._0115_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4430_  (.A(\MuI._0105_ ),
    .B(\MuI._0114_ ),
    .Y(\MuI._0116_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4431_  (.A(\MuI._0115_ ),
    .B(\MuI._0116_ ),
    .X(\MuI._0117_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4432_  (.A(\MuI._0094_ ),
    .B(\MuI._0095_ ),
    .C(\MuI._0117_ ),
    .Y(\MuI._0118_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4433_  (.A(\MuI._0094_ ),
    .B(\MuI._0118_ ),
    .Y(\MuI._0120_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4434_  (.A1(\MuI._0064_ ),
    .A2(\MuI._0066_ ),
    .B1(\MuI._0068_ ),
    .X(\MuI._0121_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4435_  (.A1(\MuI._3357_ ),
    .A2(\MuI._3358_ ),
    .B1(\MuI._3377_ ),
    .X(\MuI._0122_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._4436_  (.A1(\MuI._0121_ ),
    .A2(\MuI._0071_ ),
    .B1(\MuI._3378_ ),
    .C1(\MuI._0122_ ),
    .Y(\MuI._0123_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._4437_  (.A1(\MuI._3378_ ),
    .A2(\MuI._0122_ ),
    .B1(\MuI._0121_ ),
    .C1(\MuI._0071_ ),
    .X(\MuI._0124_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4438_  (.A(\MuI._0123_ ),
    .B(\MuI._0124_ ),
    .Y(\MuI._0125_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4439_  (.A(\MuI._0120_ ),
    .B(\MuI._0125_ ),
    .Y(\MuI._0126_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4440_  (.A(\MuI._0075_ ),
    .B(\MuI._0076_ ),
    .Y(\MuI._0127_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4441_  (.A1(\MuI._0077_ ),
    .A2(\MuI._0126_ ),
    .B1(\MuI._0127_ ),
    .Y(\MuI._0128_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4442_  (.A(\MuI._3390_ ),
    .B(\MuI._3421_ ),
    .X(\MuI._0129_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4443_  (.A(\MuI._0128_ ),
    .B(\MuI._0129_ ),
    .Y(\MuI._0131_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4444_  (.A1(\MuI._0120_ ),
    .A2(\MuI._0124_ ),
    .B1_N(\MuI._0123_ ),
    .X(\MuI._0132_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._4445_  (.A1(\MuI._3239_ ),
    .A2(\MuI._3359_ ),
    .A3(\MuI._3366_ ),
    .B1(\MuI._3375_ ),
    .X(\MuI._0133_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4446_  (.A(\MuI._0132_ ),
    .B(\MuI._0133_ ),
    .X(\MuI._0134_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4447_  (.A1(\MuI._3368_ ),
    .A2(\MuI._3373_ ),
    .B1_N(\MuI._3369_ ),
    .X(\MuI._0135_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4448_  (.A(\MuI._0134_ ),
    .B(\MuI._0135_ ),
    .Y(\MuI._0136_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4449_  (.A_N(\MuI._0128_ ),
    .B(\MuI._0129_ ),
    .X(\MuI._0137_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4450_  (.A1(\MuI._0131_ ),
    .A2(\MuI._0136_ ),
    .B1(\MuI._0137_ ),
    .X(\MuI._0138_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4451_  (.A(\MuI._0016_ ),
    .B_N(\MuI._0138_ ),
    .X(\MuI._0139_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4452_  (.A(\MuI._0138_ ),
    .B(\MuI._0016_ ),
    .X(\MuI._0140_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4453_  (.A(\MuI._0135_ ),
    .B_N(\MuI._0134_ ),
    .X(\MuI._0142_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4454_  (.A1(\MuI._0132_ ),
    .A2(\MuI._0133_ ),
    .B1(\MuI._0142_ ),
    .Y(\MuI._0143_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4455_  (.A(\MuI._0140_ ),
    .B_N(\MuI._0143_ ),
    .X(\MuI._0144_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4456_  (.A(\MuI._0015_ ),
    .B(\MuI._0139_ ),
    .C(\MuI._0144_ ),
    .X(\MuI._0145_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4457_  (.A1(\MuI._0139_ ),
    .A2(\MuI._0144_ ),
    .B1(\MuI._0015_ ),
    .Y(\MuI._0146_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4458_  (.A(\MuI._0145_ ),
    .B(\MuI._0146_ ),
    .X(\MuI._0147_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4459_  (.A(\MuI._0143_ ),
    .B(\MuI._0140_ ),
    .X(\MuI._0148_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4460_  (.A1(\MuI.a_operand[20] ),
    .A2(\MuI.b_operand[1] ),
    .B1(\MuI.b_operand[0] ),
    .B2(\MuI.a_operand[21] ),
    .X(\MuI._0149_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4461_  (.A(\MuI.a_operand[21] ),
    .B(\MuI.a_operand[20] ),
    .C(\MuI.b_operand[1] ),
    .D(\MuI.b_operand[0] ),
    .X(\MuI._0150_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4462_  (.A1(\MuI._1021_ ),
    .A2(\MuI._3269_ ),
    .A3(\MuI._0149_ ),
    .B1(\MuI._0150_ ),
    .X(\MuI._0151_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4463_  (.A1_N(\MuI._0768_ ),
    .A2_N(\MuI._3268_ ),
    .B1(\MuI._0019_ ),
    .B2(\MuI._0022_ ),
    .X(\MuI._0153_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4464_  (.A(\MuI._0023_ ),
    .B(\MuI._0153_ ),
    .Y(\MuI._0154_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4465_  (.A(\MuI._0151_ ),
    .B(\MuI._0154_ ),
    .Y(\MuI._0155_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4466_  (.A(\MuI._2066_ ),
    .B(\MuI._2895_ ),
    .Y(\MuI._0156_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4467_  (.A1(\MuI._1461_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI.a_operand[19] ),
    .Y(\MuI._0157_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4468_  (.A(\MuI.a_operand[19] ),
    .B(\MuI.a_operand[18] ),
    .C(\MuI._2884_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._0158_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4469_  (.A(\MuI._0157_ ),
    .B(\MuI._0158_ ),
    .X(\MuI._0159_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4470_  (.A(\MuI._0156_ ),
    .B(\MuI._0159_ ),
    .Y(\MuI._0160_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4471_  (.A(\MuI._0156_ ),
    .B(\MuI._0159_ ),
    .X(\MuI._0161_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4472_  (.A(\MuI._0151_ ),
    .B(\MuI._0154_ ),
    .Y(\MuI._0162_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._4473_  (.A1(\MuI._0155_ ),
    .A2(\MuI._0160_ ),
    .A3(\MuI._0161_ ),
    .B1(\MuI._0162_ ),
    .X(\MuI._0164_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4474_  (.A(\MuI._0024_ ),
    .B(\MuI._0026_ ),
    .Y(\MuI._0165_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4475_  (.A(\MuI._0165_ ),
    .B(\MuI._0033_ ),
    .Y(\MuI._0166_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4476_  (.A(\MuI._0164_ ),
    .B(\MuI._0166_ ),
    .Y(\MuI._0167_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4477_  (.A(\MuI.b_operand[8] ),
    .X(\MuI._0168_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4478_  (.A(\MuI._2671_ ),
    .B(\MuI._0168_ ),
    .Y(\MuI._0169_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4479_  (.A1(\MuI._2605_ ),
    .A2(\MuI._2873_ ),
    .B1(\MuI._2875_ ),
    .B2(\MuI._2852_ ),
    .Y(\MuI._0170_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4480_  (.A(\MuI._2852_ ),
    .B(\MuI._2605_ ),
    .C(\MuI._3189_ ),
    .D(\MuI._2868_ ),
    .X(\MuI._0171_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4481_  (.A1(\MuI._0169_ ),
    .A2(\MuI._0170_ ),
    .B1_N(\MuI._0171_ ),
    .X(\MuI._0172_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4482_  (.A(\MuI._0040_ ),
    .B(\MuI._0039_ ),
    .Y(\MuI._0173_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4483_  (.A(\MuI._0038_ ),
    .B(\MuI._0173_ ),
    .Y(\MuI._0175_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4484_  (.A1(\MuI._0158_ ),
    .A2(\MuI._0160_ ),
    .B1(\MuI._0175_ ),
    .Y(\MuI._0176_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4485_  (.A(\MuI._0158_ ),
    .B(\MuI._0160_ ),
    .C(\MuI._0175_ ),
    .X(\MuI._0177_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4486_  (.A(\MuI._0176_ ),
    .B(\MuI._0177_ ),
    .X(\MuI._0178_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4487_  (.A(\MuI._0172_ ),
    .B(\MuI._0178_ ),
    .Y(\MuI._0179_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4488_  (.A(\MuI._0164_ ),
    .B_N(\MuI._0166_ ),
    .X(\MuI._0180_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4489_  (.A1(\MuI._0167_ ),
    .A2(\MuI._0179_ ),
    .B1_N(\MuI._0180_ ),
    .Y(\MuI._0181_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4490_  (.A(\MuI._0037_ ),
    .B(\MuI._0047_ ),
    .Y(\MuI._0182_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4491_  (.A(\MuI._0181_ ),
    .B(\MuI._0182_ ),
    .X(\MuI._0183_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4492_  (.A(\MuI._2850_ ),
    .B(\MuI._2495_ ),
    .Y(\MuI._0184_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4493_  (.A1(\MuI._2975_ ),
    .A2(\MuI._2451_ ),
    .B1(\MuI._2845_ ),
    .B2(\MuI._2440_ ),
    .Y(\MuI._0186_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4494_  (.A(\MuI._2440_ ),
    .B(\MuI._2844_ ),
    .C(\MuI._2451_ ),
    .D(\MuI._2845_ ),
    .X(\MuI._0187_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4495_  (.A1(\MuI._0184_ ),
    .A2(\MuI._0186_ ),
    .B1_N(\MuI._0187_ ),
    .X(\MuI._0188_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4496_  (.A(\MuI._0055_ ),
    .B(\MuI._0053_ ),
    .Y(\MuI._0189_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4497_  (.A(\MuI._0052_ ),
    .B(\MuI._0189_ ),
    .Y(\MuI._0190_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4498_  (.A(\MuI._0188_ ),
    .B_N(\MuI._0190_ ),
    .X(\MuI._0191_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4499_  (.A(\MuI._0190_ ),
    .B(\MuI._0188_ ),
    .Y(\MuI._0192_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4500_  (.A(\MuI._0080_ ),
    .B(\MuI._0079_ ),
    .Y(\MuI._0193_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4501_  (.A(\MuI._0078_ ),
    .B(\MuI._0193_ ),
    .Y(\MuI._0194_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4502_  (.A(\MuI._0192_ ),
    .B(\MuI._0194_ ),
    .Y(\MuI._0195_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4503_  (.A(\MuI._0172_ ),
    .B_N(\MuI._0178_ ),
    .X(\MuI._0197_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4504_  (.A(\MuI._0060_ ),
    .B(\MuI._0062_ ),
    .X(\MuI._0198_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4505_  (.A(\MuI._0063_ ),
    .B(\MuI._0198_ ),
    .Y(\MuI._0199_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4506_  (.A1(\MuI._0176_ ),
    .A2(\MuI._0197_ ),
    .B1(\MuI._0199_ ),
    .Y(\MuI._0200_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4507_  (.A(\MuI._0176_ ),
    .B(\MuI._0197_ ),
    .C(\MuI._0199_ ),
    .X(\MuI._0201_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4508_  (.A1(\MuI._0191_ ),
    .A2(\MuI._0195_ ),
    .B1(\MuI._0200_ ),
    .C1(\MuI._0201_ ),
    .X(\MuI._0202_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4509_  (.A1(\MuI._0200_ ),
    .A2(\MuI._0201_ ),
    .B1(\MuI._0191_ ),
    .C1(\MuI._0195_ ),
    .Y(\MuI._0203_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4510_  (.A(\MuI._0202_ ),
    .B(\MuI._0203_ ),
    .X(\MuI._0204_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4511_  (.A(\MuI._0181_ ),
    .B(\MuI._0182_ ),
    .Y(\MuI._0205_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4512_  (.A1(\MuI._0183_ ),
    .A2(\MuI._0204_ ),
    .B1(\MuI._0205_ ),
    .X(\MuI._0206_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4513_  (.A(\MuI._0051_ ),
    .B(\MuI._0073_ ),
    .X(\MuI._0208_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4514_  (.A(\MuI._0206_ ),
    .B(\MuI._0208_ ),
    .X(\MuI._0209_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4515_  (.A(\MuI.b_operand[14] ),
    .B(\MuI._2352_ ),
    .Y(\MuI._0210_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._4516_  (.A1(\MuI._2649_ ),
    .A2(\MuI._2773_ ),
    .B1(\MuI._2786_ ),
    .B2(\MuI._2704_ ),
    .Y(\MuI._0211_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4517_  (.A(\MuI._2799_ ),
    .B(\MuI._2918_ ),
    .C(\MuI._2790_ ),
    .D(\MuI._3223_ ),
    .X(\MuI._0212_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4518_  (.A1(\MuI._0210_ ),
    .A2(\MuI._0211_ ),
    .B1_N(\MuI._0212_ ),
    .X(\MuI._0213_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4519_  (.A1_N(\MuI._1263_ ),
    .A2_N(\MuI._3363_ ),
    .B1(\MuI._0087_ ),
    .B2(\MuI._0089_ ),
    .X(\MuI._0214_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4520_  (.A(\MuI._0213_ ),
    .B(\MuI._0090_ ),
    .C(\MuI._0214_ ),
    .X(\MuI._0215_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4521_  (.A(\MuI._3000_ ),
    .B(\MuI._1791_ ),
    .C(\MuI._0088_ ),
    .D(\MuI._3362_ ),
    .X(\MuI._0216_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4522_  (.A1(\MuI._1802_ ),
    .A2(\MuI._2374_ ),
    .B1(\MuI._3363_ ),
    .B2(\MuI._1307_ ),
    .Y(\MuI._0217_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4523_  (.A_N(\MuI._0216_ ),
    .B_N(\MuI._0217_ ),
    .C(\MuI._1263_ ),
    .D(\MuI._0101_ ),
    .X(\MuI._0219_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4524_  (.A(\MuI._0216_ ),
    .B(\MuI._0219_ ),
    .X(\MuI._0220_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4525_  (.A(\MuI._0090_ ),
    .B(\MuI._0214_ ),
    .Y(\MuI._0221_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4526_  (.A(\MuI._0213_ ),
    .B(\MuI._0221_ ),
    .Y(\MuI._0222_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4527_  (.A(\MuI._0220_ ),
    .B(\MuI._0222_ ),
    .Y(\MuI._0223_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4528_  (.A(\MuI._0087_ ),
    .B(\MuI._0090_ ),
    .C(\MuI._0091_ ),
    .X(\MuI._0224_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4529_  (.A(\MuI._0092_ ),
    .B(\MuI._0224_ ),
    .Y(\MuI._0225_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4530_  (.A1(\MuI._0215_ ),
    .A2(\MuI._0223_ ),
    .B1(\MuI._0225_ ),
    .Y(\MuI._0226_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4531_  (.A(\MuI._0215_ ),
    .B(\MuI._0223_ ),
    .C(\MuI._0225_ ),
    .X(\MuI._0227_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4532_  (.A(\MuI.a_operand[4] ),
    .X(\MuI._0228_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4533_  (.A(\MuI.b_operand[19] ),
    .B(\MuI._2811_ ),
    .C(\MuI._2829_ ),
    .D(\MuI._0228_ ),
    .X(\MuI._0230_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4534_  (.A1(\MuI._1142_ ),
    .A2(\MuI._0101_ ),
    .B1(\MuI._3246_ ),
    .B2(\MuI._2939_ ),
    .Y(\MuI._0231_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4535_  (.A(\MuI._0230_ ),
    .B(\MuI._0231_ ),
    .Y(\MuI._0232_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4536_  (.A(\MuI._2817_ ),
    .B(\MuI._3372_ ),
    .C(\MuI._0232_ ),
    .X(\MuI._0233_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4537_  (.A(\MuI._0103_ ),
    .B(\MuI._0102_ ),
    .Y(\MuI._0234_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4538_  (.A(\MuI._0099_ ),
    .B(\MuI._0234_ ),
    .Y(\MuI._0235_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4539_  (.A1(\MuI._0230_ ),
    .A2(\MuI._0233_ ),
    .B1(\MuI._0235_ ),
    .X(\MuI._0236_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4540_  (.A(\MuI._0230_ ),
    .B(\MuI._0233_ ),
    .C(\MuI._0235_ ),
    .Y(\MuI._0237_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4541_  (.A(\MuI._0236_ ),
    .B(\MuI._0237_ ),
    .Y(\MuI._0238_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4542_  (.A1(\MuI.b_operand[21] ),
    .A2(\MuI._3372_ ),
    .B1(\MuI._0111_ ),
    .B2(\MuI.b_operand[22] ),
    .X(\MuI._0239_ ));
 sky130_fd_sc_hd__inv_2 \MuI._4543_  (.A(\MuI._0239_ ),
    .Y(\MuI._0241_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4544_  (.A(\MuI._2826_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._3372_ ),
    .D(\MuI._0112_ ),
    .X(\MuI._0242_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4545_  (.A(\MuI._0241_ ),
    .B(\MuI._0242_ ),
    .Y(\MuI._0243_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4546_  (.A(\MuI.a_operand[1] ),
    .X(\MuI._0244_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4547_  (.A(\MuI._0244_ ),
    .X(\MuI._0245_ ));
 sky130_fd_sc_hd__buf_4 \MuI._4548_  (.A(\MuI._0245_ ),
    .X(\MuI._0246_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4549_  (.A(\MuI._0246_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._0247_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4550_  (.A(\MuI._0243_ ),
    .B(\MuI._0247_ ),
    .Y(\MuI._0248_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4551_  (.A(\MuI._0238_ ),
    .B(\MuI._0248_ ),
    .X(\MuI._0249_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4552_  (.A(\MuI._0238_ ),
    .B(\MuI._0248_ ),
    .Y(\MuI._0250_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4553_  (.A(\MuI._0249_ ),
    .B(\MuI._0250_ ),
    .X(\MuI._0252_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4554_  (.A(\MuI._0226_ ),
    .B(\MuI._0227_ ),
    .C(\MuI._0252_ ),
    .Y(\MuI._0253_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4555_  (.A(\MuI._0226_ ),
    .B(\MuI._0253_ ),
    .X(\MuI._0254_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4556_  (.A1(\MuI._0176_ ),
    .A2(\MuI._0197_ ),
    .B1(\MuI._0199_ ),
    .X(\MuI._0255_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4557_  (.A1(\MuI._0094_ ),
    .A2(\MuI._0095_ ),
    .B1(\MuI._0117_ ),
    .X(\MuI._0256_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4558_  (.A(\MuI._0118_ ),
    .B(\MuI._0256_ ),
    .X(\MuI._0257_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4559_  (.A1(\MuI._0255_ ),
    .A2(\MuI._0202_ ),
    .B1(\MuI._0257_ ),
    .Y(\MuI._0258_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4560_  (.A(\MuI._0255_ ),
    .B(\MuI._0202_ ),
    .C(\MuI._0257_ ),
    .X(\MuI._0259_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4561_  (.A(\MuI._0258_ ),
    .B(\MuI._0259_ ),
    .Y(\MuI._0260_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4562_  (.A(\MuI._0254_ ),
    .B(\MuI._0260_ ),
    .X(\MuI._0261_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4563_  (.A(\MuI._0206_ ),
    .B(\MuI._0208_ ),
    .Y(\MuI._0263_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4564_  (.A1(\MuI._0209_ ),
    .A2(\MuI._0261_ ),
    .B1_N(\MuI._0263_ ),
    .Y(\MuI._0264_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4565_  (.A(\MuI._0077_ ),
    .B(\MuI._0126_ ),
    .X(\MuI._0265_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4566_  (.A(\MuI._0264_ ),
    .B(\MuI._0265_ ),
    .Y(\MuI._0266_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4567_  (.A1(\MuI._0254_ ),
    .A2(\MuI._0260_ ),
    .B1(\MuI._0258_ ),
    .X(\MuI._0267_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4568_  (.A_N(\MuI._0104_ ),
    .B(\MuI._0098_ ),
    .X(\MuI._0268_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4569_  (.A(\MuI._0268_ ),
    .B(\MuI._0115_ ),
    .Y(\MuI._0269_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4570_  (.A(\MuI._0267_ ),
    .B(\MuI._0269_ ),
    .Y(\MuI._0270_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4571_  (.A1(\MuI._0112_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._0109_ ),
    .B1(\MuI._0107_ ),
    .X(\MuI._0271_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4572_  (.A(\MuI._0270_ ),
    .B(\MuI._0271_ ),
    .X(\MuI._0272_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4573_  (.A_N(\MuI._0264_ ),
    .B(\MuI._0265_ ),
    .X(\MuI._0274_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4574_  (.A1(\MuI._0266_ ),
    .A2(\MuI._0272_ ),
    .B1(\MuI._0274_ ),
    .X(\MuI._0275_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4575_  (.A(\MuI._0131_ ),
    .B(\MuI._0136_ ),
    .X(\MuI._0276_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4576_  (.A(\MuI._0275_ ),
    .B(\MuI._0276_ ),
    .Y(\MuI._0277_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4577_  (.A1(\MuI._0268_ ),
    .A2(\MuI._0115_ ),
    .B1(\MuI._0267_ ),
    .Y(\MuI._0278_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4578_  (.A1(\MuI._0270_ ),
    .A2(\MuI._0271_ ),
    .B1_N(\MuI._0278_ ),
    .X(\MuI._0279_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4579_  (.A(\MuI._0277_ ),
    .B_N(\MuI._0279_ ),
    .X(\MuI._0280_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4580_  (.A1(\MuI._0275_ ),
    .A2(\MuI._0276_ ),
    .B1_N(\MuI._0280_ ),
    .Y(\MuI._0281_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4581_  (.A(\MuI._0148_ ),
    .B(\MuI._0281_ ),
    .Y(\MuI._0282_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4582_  (.A(\MuI._0014_ ),
    .B(\MuI._0147_ ),
    .C(\MuI._0282_ ),
    .Y(\MuI._0283_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4583_  (.A(\MuI._0279_ ),
    .B(\MuI._0277_ ),
    .X(\MuI._0285_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4584_  (.A(\MuI._2796_ ),
    .B(\MuI._2374_ ),
    .Y(\MuI._0286_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4585_  (.A1(\MuI._2803_ ),
    .A2(\MuI._2786_ ),
    .B1(\MuI._2352_ ),
    .B2(\MuI._2802_ ),
    .Y(\MuI._0287_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4586_  (.A(\MuI._2799_ ),
    .B(\MuI._2918_ ),
    .C(\MuI._3223_ ),
    .D(\MuI._3349_ ),
    .X(\MuI._0288_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4587_  (.A1(\MuI._0286_ ),
    .A2(\MuI._0287_ ),
    .B1_N(\MuI._0288_ ),
    .X(\MuI._0289_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4588_  (.A1_N(\MuI._2473_ ),
    .A2_N(\MuI._2830_ ),
    .B1(\MuI._0216_ ),
    .B2(\MuI._0217_ ),
    .X(\MuI._0290_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4589_  (.A(\MuI._0219_ ),
    .B(\MuI._0289_ ),
    .C(\MuI._0290_ ),
    .X(\MuI._0291_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4590_  (.A(\MuI._1296_ ),
    .B(\MuI._1791_ ),
    .C(\MuI._3362_ ),
    .D(\MuI._2829_ ),
    .X(\MuI._0292_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4591_  (.A1(\MuI._1802_ ),
    .A2(\MuI._2319_ ),
    .B1(\MuI._0101_ ),
    .B2(\MuI._1307_ ),
    .Y(\MuI._0293_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4592_  (.A_N(\MuI._0292_ ),
    .B_N(\MuI._0293_ ),
    .C(\MuI._1263_ ),
    .D(\MuI._3246_ ),
    .X(\MuI._0294_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4593_  (.A(\MuI._0292_ ),
    .B(\MuI._0294_ ),
    .X(\MuI._0296_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4594_  (.A(\MuI._0219_ ),
    .B(\MuI._0290_ ),
    .Y(\MuI._0297_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4595_  (.A(\MuI._0289_ ),
    .B(\MuI._0297_ ),
    .Y(\MuI._0298_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4596_  (.A(\MuI._0296_ ),
    .B(\MuI._0298_ ),
    .Y(\MuI._0299_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4597_  (.A(\MuI._0220_ ),
    .B(\MuI._0222_ ),
    .Y(\MuI._0300_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4598_  (.A1(\MuI._0291_ ),
    .A2(\MuI._0299_ ),
    .B1(\MuI._0300_ ),
    .Y(\MuI._0301_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4599_  (.A(\MuI._0300_ ),
    .B(\MuI._0291_ ),
    .C(\MuI._0299_ ),
    .X(\MuI._0302_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4600_  (.A(\MuI.b_operand[19] ),
    .B(\MuI.b_operand[18] ),
    .C(\MuI._0228_ ),
    .D(\MuI._3371_ ),
    .X(\MuI._0303_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4601_  (.A(\MuI.a_operand[3] ),
    .X(\MuI._0304_ ));
 sky130_fd_sc_hd__buf_4 \MuI._4602_  (.A(\MuI._0304_ ),
    .X(\MuI._0305_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4603_  (.A1(\MuI._2811_ ),
    .A2(\MuI._3246_ ),
    .B1(\MuI._0305_ ),
    .B2(\MuI._2939_ ),
    .Y(\MuI._0307_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4604_  (.A(\MuI._0303_ ),
    .B(\MuI._0307_ ),
    .Y(\MuI._0308_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4605_  (.A(\MuI._0867_ ),
    .B(\MuI._0111_ ),
    .C(\MuI._0308_ ),
    .X(\MuI._0309_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4606_  (.A(\MuI.b_operand[20] ),
    .B(\MuI._3372_ ),
    .Y(\MuI._0310_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4607_  (.A(\MuI._0232_ ),
    .B(\MuI._0310_ ),
    .Y(\MuI._0311_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4608_  (.A1(\MuI._0303_ ),
    .A2(\MuI._0309_ ),
    .B1(\MuI._0311_ ),
    .X(\MuI._0312_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4609_  (.A(\MuI._0311_ ),
    .B(\MuI._0303_ ),
    .C(\MuI._0309_ ),
    .Y(\MuI._0313_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4610_  (.A(\MuI._0312_ ),
    .B(\MuI._0313_ ),
    .Y(\MuI._0314_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4611_  (.A(\MuI._0244_ ),
    .X(\MuI._0315_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4612_  (.A(\MuI._2826_ ),
    .B(\MuI.b_operand[21] ),
    .C(\MuI._0315_ ),
    .X(\MuI._0316_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4613_  (.A1(\MuI.b_operand[21] ),
    .A2(\MuI._0111_ ),
    .B1(\MuI._0315_ ),
    .B2(\MuI._2826_ ),
    .X(\MuI._0318_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4614_  (.A1(\MuI._0112_ ),
    .A2(\MuI._0316_ ),
    .B1_N(\MuI._0318_ ),
    .X(\MuI._0319_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4615_  (.A(\MuI.a_operand[0] ),
    .X(\MuI._0320_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4616_  (.A(\MuI._0320_ ),
    .X(\MuI._0321_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4617_  (.A(\MuI._0321_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._0322_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4618_  (.A(\MuI._0319_ ),
    .B(\MuI._0322_ ),
    .Y(\MuI._0323_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4619_  (.A(\MuI._0314_ ),
    .B(\MuI._0323_ ),
    .X(\MuI._0324_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4620_  (.A(\MuI._0301_ ),
    .B(\MuI._0302_ ),
    .C(\MuI._0324_ ),
    .Y(\MuI._0325_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4621_  (.A(\MuI._0301_ ),
    .B(\MuI._0325_ ),
    .X(\MuI._0326_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4622_  (.A(\MuI.a_operand[12] ),
    .X(\MuI._0327_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4623_  (.A(\MuI.b_operand[10] ),
    .B(\MuI._0327_ ),
    .C(\MuI._2837_ ),
    .D(\MuI.a_operand[11] ),
    .X(\MuI._0329_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4624_  (.A1(\MuI._0327_ ),
    .A2(\MuI._2854_ ),
    .B1(\MuI._2484_ ),
    .B2(\MuI._2853_ ),
    .Y(\MuI._0330_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4625_  (.A_N(\MuI._0329_ ),
    .B_N(\MuI._0330_ ),
    .C(\MuI.b_operand[11] ),
    .D(\MuI._2790_ ),
    .X(\MuI._0331_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4626_  (.A(\MuI._0329_ ),
    .B(\MuI._0331_ ),
    .Y(\MuI._0332_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4627_  (.A(\MuI._0187_ ),
    .B(\MuI._0186_ ),
    .Y(\MuI._0333_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4628_  (.A(\MuI._0184_ ),
    .B(\MuI._0333_ ),
    .Y(\MuI._0334_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4629_  (.A(\MuI._0332_ ),
    .B_N(\MuI._0334_ ),
    .X(\MuI._0335_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4630_  (.A(\MuI._0334_ ),
    .B(\MuI._0332_ ),
    .Y(\MuI._0336_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4631_  (.A(\MuI._0212_ ),
    .B(\MuI._0211_ ),
    .Y(\MuI._0337_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4632_  (.A(\MuI._0210_ ),
    .B(\MuI._0337_ ),
    .Y(\MuI._0338_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4633_  (.A(\MuI._0336_ ),
    .B(\MuI._0338_ ),
    .Y(\MuI._0340_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4634_  (.A(\MuI._0335_ ),
    .B(\MuI._0340_ ),
    .Y(\MuI._0341_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4635_  (.A(\MuI.a_operand[18] ),
    .B(\MuI.a_operand[17] ),
    .C(\MuI._2884_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._0342_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4636_  (.A(\MuI._2840_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._0343_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4637_  (.A1(\MuI.a_operand[17] ),
    .A2(\MuI._2884_ ),
    .B1(\MuI._3307_ ),
    .B2(\MuI._1461_ ),
    .Y(\MuI._0344_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4638_  (.A(\MuI._0344_ ),
    .B(\MuI._0342_ ),
    .X(\MuI._0345_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4639_  (.A(\MuI._0343_ ),
    .B(\MuI._0345_ ),
    .Y(\MuI._0346_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4640_  (.A(\MuI._0171_ ),
    .B(\MuI._0170_ ),
    .Y(\MuI._0347_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4641_  (.A(\MuI._0169_ ),
    .B(\MuI._0347_ ),
    .Y(\MuI._0348_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4642_  (.A1(\MuI._0342_ ),
    .A2(\MuI._0346_ ),
    .B1(\MuI._0348_ ),
    .Y(\MuI._0349_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4643_  (.A(\MuI._2440_ ),
    .B(\MuI.b_operand[8] ),
    .Y(\MuI._0351_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4644_  (.A1(\MuI.a_operand[14] ),
    .A2(\MuI._2866_ ),
    .B1(\MuI._2868_ ),
    .B2(\MuI.a_operand[15] ),
    .Y(\MuI._0352_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4645_  (.A(\MuI.a_operand[15] ),
    .B(\MuI.a_operand[14] ),
    .C(\MuI._2866_ ),
    .D(\MuI.b_operand[6] ),
    .X(\MuI._0353_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._4646_  (.A1(\MuI._0351_ ),
    .A2(\MuI._0352_ ),
    .B1_N(\MuI._0353_ ),
    .X(\MuI._0354_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4647_  (.A(\MuI._0342_ ),
    .B(\MuI._0346_ ),
    .C(\MuI._0348_ ),
    .X(\MuI._0355_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4648_  (.A(\MuI._0349_ ),
    .B(\MuI._0355_ ),
    .X(\MuI._0356_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4649_  (.A(\MuI._0354_ ),
    .B_N(\MuI._0356_ ),
    .X(\MuI._0357_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4650_  (.A(\MuI._0192_ ),
    .B(\MuI._0194_ ),
    .X(\MuI._0358_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4651_  (.A(\MuI._0195_ ),
    .B(\MuI._0358_ ),
    .Y(\MuI._0359_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4652_  (.A1(\MuI._0349_ ),
    .A2(\MuI._0357_ ),
    .B1(\MuI._0359_ ),
    .Y(\MuI._0360_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4653_  (.A(\MuI._0349_ ),
    .B(\MuI._0357_ ),
    .C(\MuI._0359_ ),
    .X(\MuI._0362_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4654_  (.A(\MuI._0360_ ),
    .B(\MuI._0362_ ),
    .Y(\MuI._0363_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4655_  (.A1(\MuI._0341_ ),
    .A2(\MuI._0363_ ),
    .B1(\MuI._0360_ ),
    .X(\MuI._0364_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4656_  (.A1(\MuI._0226_ ),
    .A2(\MuI._0227_ ),
    .B1(\MuI._0252_ ),
    .X(\MuI._0365_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4657_  (.A(\MuI._0253_ ),
    .B(\MuI._0365_ ),
    .X(\MuI._0366_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4658_  (.A(\MuI._0364_ ),
    .B(\MuI._0366_ ),
    .Y(\MuI._0367_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4659_  (.A_N(\MuI._0366_ ),
    .B(\MuI._0364_ ),
    .X(\MuI._0368_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4660_  (.A1(\MuI._0326_ ),
    .A2(\MuI._0367_ ),
    .B1(\MuI._0368_ ),
    .X(\MuI._0369_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4661_  (.A(\MuI._0236_ ),
    .B(\MuI._0249_ ),
    .Y(\MuI._0370_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4662_  (.A(\MuI._0369_ ),
    .B(\MuI._0370_ ),
    .Y(\MuI._0371_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4663_  (.A1(\MuI._0246_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._0239_ ),
    .B1(\MuI._0242_ ),
    .X(\MuI._0373_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4664_  (.A1(\MuI._0236_ ),
    .A2(\MuI._0249_ ),
    .B1(\MuI._0369_ ),
    .Y(\MuI._0374_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4665_  (.A1(\MuI._0371_ ),
    .A2(\MuI._0373_ ),
    .B1_N(\MuI._0374_ ),
    .X(\MuI._0375_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4666_  (.A(\MuI.a_operand[20] ),
    .B(\MuI.a_operand[19] ),
    .C(\MuI.b_operand[1] ),
    .D(\MuI.b_operand[0] ),
    .X(\MuI._0376_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4667_  (.A1(\MuI.a_operand[19] ),
    .A2(\MuI._0017_ ),
    .B1(\MuI._0018_ ),
    .B2(\MuI.a_operand[20] ),
    .Y(\MuI._0377_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4668_  (.A(\MuI.b_operand[2] ),
    .X(\MuI._0378_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4669_  (.A_N(\MuI._0376_ ),
    .B_N(\MuI._0377_ ),
    .C(\MuI._1461_ ),
    .D(\MuI._0378_ ),
    .X(\MuI._0379_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4670_  (.A(\MuI._0376_ ),
    .B(\MuI._0379_ ),
    .Y(\MuI._0380_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4671_  (.A(\MuI._1010_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._0381_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4672_  (.A_N(\MuI._0150_ ),
    .B(\MuI._0149_ ),
    .X(\MuI._0382_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4673_  (.A(\MuI._0381_ ),
    .B(\MuI._0382_ ),
    .Y(\MuI._0384_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4674_  (.A_N(\MuI._0380_ ),
    .B(\MuI._0384_ ),
    .X(\MuI._0385_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4675_  (.A(\MuI._0380_ ),
    .B(\MuI._0384_ ),
    .Y(\MuI._0386_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4676_  (.A(\MuI._0343_ ),
    .B(\MuI._0345_ ),
    .X(\MuI._0387_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4677_  (.A(\MuI._0346_ ),
    .B(\MuI._0387_ ),
    .Y(\MuI._0388_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4678_  (.A(\MuI._0386_ ),
    .B(\MuI._0388_ ),
    .X(\MuI._0389_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4679_  (.A(\MuI._0160_ ),
    .B(\MuI._0161_ ),
    .Y(\MuI._0390_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4680_  (.A(\MuI._0155_ ),
    .B(\MuI._0390_ ),
    .Y(\MuI._0391_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4681_  (.A(\MuI._0385_ ),
    .B(\MuI._0389_ ),
    .C(\MuI._0391_ ),
    .X(\MuI._0392_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4682_  (.A(\MuI._0354_ ),
    .B(\MuI._0356_ ),
    .Y(\MuI._0393_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4683_  (.A1(\MuI._0385_ ),
    .A2(\MuI._0389_ ),
    .B1(\MuI._0391_ ),
    .Y(\MuI._0395_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4684_  (.A1(\MuI._0392_ ),
    .A2(\MuI._0393_ ),
    .B1_N(\MuI._0395_ ),
    .X(\MuI._0396_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4685_  (.A(\MuI._0167_ ),
    .B(\MuI._0179_ ),
    .Y(\MuI._0397_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4686_  (.A(\MuI._0396_ ),
    .B_N(\MuI._0397_ ),
    .X(\MuI._0398_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4687_  (.A(\MuI._0341_ ),
    .B(\MuI._0363_ ),
    .X(\MuI._0399_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4688_  (.A_N(\MuI._0397_ ),
    .B(\MuI._0396_ ),
    .X(\MuI._0400_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4689_  (.A1(\MuI._0398_ ),
    .A2(\MuI._0399_ ),
    .B1(\MuI._0400_ ),
    .Y(\MuI._0401_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4690_  (.A(\MuI._0183_ ),
    .B(\MuI._0204_ ),
    .Y(\MuI._0402_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4691_  (.A(\MuI._0401_ ),
    .B(\MuI._0402_ ),
    .X(\MuI._0403_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4692_  (.A(\MuI._0326_ ),
    .B(\MuI._0367_ ),
    .X(\MuI._0404_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4693_  (.A(\MuI._0401_ ),
    .B(\MuI._0402_ ),
    .Y(\MuI._0406_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4694_  (.A1(\MuI._0403_ ),
    .A2(\MuI._0404_ ),
    .B1(\MuI._0406_ ),
    .Y(\MuI._0407_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4695_  (.A(\MuI._0209_ ),
    .B(\MuI._0261_ ),
    .X(\MuI._0408_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4696_  (.A(\MuI._0407_ ),
    .B(\MuI._0408_ ),
    .Y(\MuI._0409_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4697_  (.A(\MuI._0371_ ),
    .B(\MuI._0373_ ),
    .X(\MuI._0410_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4698_  (.A_N(\MuI._0407_ ),
    .B(\MuI._0408_ ),
    .X(\MuI._0411_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4699_  (.A1(\MuI._0409_ ),
    .A2(\MuI._0410_ ),
    .B1(\MuI._0411_ ),
    .Y(\MuI._0412_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4700_  (.A(\MuI._0266_ ),
    .B(\MuI._0272_ ),
    .Y(\MuI._0413_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4701_  (.A(\MuI._0412_ ),
    .B(\MuI._0413_ ),
    .X(\MuI._0414_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4702_  (.A(\MuI._0412_ ),
    .B(\MuI._0413_ ),
    .Y(\MuI._0415_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4703_  (.A1(\MuI._0375_ ),
    .A2(\MuI._0414_ ),
    .B1(\MuI._0415_ ),
    .Y(\MuI._0417_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4704_  (.A(\MuI._0285_ ),
    .B(\MuI._0417_ ),
    .Y(\MuI._0418_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4705_  (.A(\MuI._0375_ ),
    .B(\MuI._0414_ ),
    .Y(\MuI._0419_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4706_  (.A(\MuI._0321_ ),
    .X(\MuI._0420_ ));
 sky130_fd_sc_hd__buf_4 \MuI._4707_  (.A(\MuI._0420_ ),
    .X(\MuI._0421_ ));
 sky130_fd_sc_hd__a32o_1 \MuI._4708_  (.A1(\MuI._0421_ ),
    .A2(\MuI._0471_ ),
    .A3(\MuI._0318_ ),
    .B1(\MuI._0316_ ),
    .B2(\MuI._0112_ ),
    .X(\MuI._0422_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4709_  (.A(\MuI._2693_ ),
    .B(\MuI._2638_ ),
    .C(\MuI._3349_ ),
    .D(\MuI._0088_ ),
    .X(\MuI._0423_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4710_  (.A1(\MuI._2803_ ),
    .A2(\MuI._2352_ ),
    .B1(\MuI._2374_ ),
    .B2(\MuI._2802_ ),
    .Y(\MuI._0424_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4711_  (.A_N(\MuI._0423_ ),
    .B_N(\MuI._0424_ ),
    .C(\MuI.b_operand[14] ),
    .D(\MuI._3363_ ),
    .X(\MuI._0425_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4712_  (.A(\MuI._0423_ ),
    .B(\MuI._0425_ ),
    .Y(\MuI._0426_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4713_  (.A1_N(\MuI._2473_ ),
    .A2_N(\MuI._3247_ ),
    .B1(\MuI._0292_ ),
    .B2(\MuI._0293_ ),
    .X(\MuI._0428_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4714_  (.A(\MuI._0294_ ),
    .B(\MuI._0426_ ),
    .C(\MuI._0428_ ),
    .X(\MuI._0429_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4715_  (.A(\MuI._3000_ ),
    .B(\MuI._2754_ ),
    .C(\MuI._2829_ ),
    .D(\MuI._0228_ ),
    .X(\MuI._0430_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4716_  (.A1(\MuI._1802_ ),
    .A2(\MuI._0101_ ),
    .B1(\MuI._3246_ ),
    .B2(\MuI._2550_ ),
    .Y(\MuI._0431_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4717_  (.A_N(\MuI._0430_ ),
    .B_N(\MuI._0431_ ),
    .C(\MuI._2473_ ),
    .D(\MuI._3372_ ),
    .X(\MuI._0432_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4718_  (.A(\MuI._0430_ ),
    .B(\MuI._0432_ ),
    .X(\MuI._0433_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4719_  (.A(\MuI._0294_ ),
    .B(\MuI._0428_ ),
    .Y(\MuI._0434_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4720_  (.A(\MuI._0426_ ),
    .B(\MuI._0434_ ),
    .Y(\MuI._0435_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4721_  (.A(\MuI._0433_ ),
    .B(\MuI._0435_ ),
    .Y(\MuI._0436_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4722_  (.A(\MuI._0296_ ),
    .B(\MuI._0298_ ),
    .Y(\MuI._0437_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4723_  (.A1(\MuI._0429_ ),
    .A2(\MuI._0436_ ),
    .B1(\MuI._0437_ ),
    .Y(\MuI._0439_ ));
 sky130_fd_sc_hd__inv_2 \MuI._4724_  (.A(\MuI._0439_ ),
    .Y(\MuI._0440_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4725_  (.A(\MuI._0437_ ),
    .B(\MuI._0429_ ),
    .C(\MuI._0436_ ),
    .Y(\MuI._0441_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4726_  (.A1(\MuI._0878_ ),
    .A2(\MuI._0112_ ),
    .B1(\MuI._0308_ ),
    .Y(\MuI._0442_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4727_  (.A(\MuI._0309_ ),
    .B(\MuI._0442_ ),
    .X(\MuI._0443_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4728_  (.A(\MuI.a_operand[2] ),
    .X(\MuI._0444_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._4729_  (.A(\MuI._0444_ ),
    .X(\MuI._0445_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4730_  (.A1(\MuI._1142_ ),
    .A2(\MuI._0305_ ),
    .B1(\MuI._0445_ ),
    .B2(\MuI._2939_ ),
    .X(\MuI._0446_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4731_  (.A(\MuI._2939_ ),
    .B(\MuI._1142_ ),
    .C(\MuI._0305_ ),
    .D(\MuI._0445_ ),
    .X(\MuI._0447_ ));
 sky130_fd_sc_hd__a31oi_2 \MuI._4732_  (.A1(\MuI._0878_ ),
    .A2(\MuI._0246_ ),
    .A3(\MuI._0446_ ),
    .B1(\MuI._0447_ ),
    .Y(\MuI._0448_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4733_  (.A(\MuI._0443_ ),
    .B(\MuI._0448_ ),
    .Y(\MuI._0450_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4734_  (.A1(\MuI._0625_ ),
    .A2(\MuI._0246_ ),
    .B1(\MuI._0420_ ),
    .B2(\MuI._0372_ ),
    .Y(\MuI._0451_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4735_  (.A(\MuI._0321_ ),
    .B(\MuI._0316_ ),
    .X(\MuI._0452_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4736_  (.A(\MuI._0451_ ),
    .B(\MuI._0452_ ),
    .X(\MuI._0453_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4737_  (.A(\MuI._0450_ ),
    .B(\MuI._0453_ ),
    .X(\MuI._0454_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4738_  (.A(\MuI._0440_ ),
    .B(\MuI._0441_ ),
    .C(\MuI._0454_ ),
    .X(\MuI._0455_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4739_  (.A(\MuI._0439_ ),
    .B(\MuI._0455_ ),
    .X(\MuI._0456_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4740_  (.A(\MuI.a_operand[17] ),
    .B(\MuI.a_operand[16] ),
    .C(\MuI.b_operand[4] ),
    .D(\MuI._2880_ ),
    .X(\MuI._0457_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4741_  (.A(\MuI._2616_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._0458_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4742_  (.A1(\MuI._2852_ ),
    .A2(\MuI._2884_ ),
    .B1(\MuI._2880_ ),
    .B2(\MuI.a_operand[17] ),
    .Y(\MuI._0459_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4743_  (.A(\MuI._0457_ ),
    .B(\MuI._0459_ ),
    .X(\MuI._0461_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4744_  (.A(\MuI._0458_ ),
    .B(\MuI._0461_ ),
    .Y(\MuI._0462_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4745_  (.A(\MuI._0353_ ),
    .B(\MuI._0352_ ),
    .Y(\MuI._0463_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4746_  (.A(\MuI._0351_ ),
    .B(\MuI._0463_ ),
    .Y(\MuI._0464_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4747_  (.A1(\MuI._0457_ ),
    .A2(\MuI._0462_ ),
    .B1(\MuI._0464_ ),
    .Y(\MuI._0465_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4748_  (.A(\MuI.a_operand[14] ),
    .B(\MuI.a_operand[13] ),
    .C(\MuI._2866_ ),
    .D(\MuI._2868_ ),
    .X(\MuI._0466_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4749_  (.A1(\MuI._2429_ ),
    .A2(\MuI._3189_ ),
    .B1(\MuI._3190_ ),
    .B2(\MuI._2660_ ),
    .Y(\MuI._0467_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4750_  (.A_N(\MuI._0466_ ),
    .B_N(\MuI._0467_ ),
    .C(\MuI._2451_ ),
    .D(\MuI.b_operand[8] ),
    .X(\MuI._0468_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4751_  (.A(\MuI._0466_ ),
    .B(\MuI._0468_ ),
    .Y(\MuI._0469_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4752_  (.A(\MuI._0457_ ),
    .B(\MuI._0462_ ),
    .C(\MuI._0464_ ),
    .X(\MuI._0470_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4753_  (.A(\MuI._0465_ ),
    .B(\MuI._0470_ ),
    .X(\MuI._0472_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4754_  (.A(\MuI._0469_ ),
    .B_N(\MuI._0472_ ),
    .X(\MuI._0473_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4755_  (.A(\MuI._0336_ ),
    .B(\MuI._0338_ ),
    .X(\MuI._0474_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4756_  (.A(\MuI._0340_ ),
    .B(\MuI._0474_ ),
    .Y(\MuI._0475_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4757_  (.A1(\MuI._0465_ ),
    .A2(\MuI._0473_ ),
    .B1(\MuI._0475_ ),
    .X(\MuI._0476_ ));
 sky130_fd_sc_hd__buf_2 \MuI._4758_  (.A(\MuI.a_operand[11] ),
    .X(\MuI._0477_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4759_  (.A(\MuI.b_operand[10] ),
    .B(\MuI._2837_ ),
    .C(\MuI._0477_ ),
    .D(\MuI.a_operand[10] ),
    .X(\MuI._0478_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4760_  (.A1(\MuI._2854_ ),
    .A2(\MuI._0477_ ),
    .B1(\MuI._2790_ ),
    .B2(\MuI._2836_ ),
    .Y(\MuI._0479_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4761_  (.A_N(\MuI._0478_ ),
    .B_N(\MuI._0479_ ),
    .C(\MuI.b_operand[11] ),
    .D(\MuI._3223_ ),
    .X(\MuI._0480_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4762_  (.A(\MuI._0478_ ),
    .B(\MuI._0480_ ),
    .Y(\MuI._0481_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4763_  (.A1_N(\MuI._2841_ ),
    .A2_N(\MuI._2773_ ),
    .B1(\MuI._0329_ ),
    .B2(\MuI._0330_ ),
    .X(\MuI._0483_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4764_  (.A(\MuI._0331_ ),
    .B(\MuI._0483_ ),
    .Y(\MuI._0484_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4765_  (.A_N(\MuI._0481_ ),
    .B(\MuI._0484_ ),
    .X(\MuI._0485_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4766_  (.A(\MuI._0484_ ),
    .B(\MuI._0481_ ),
    .Y(\MuI._0486_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4767_  (.A(\MuI._0288_ ),
    .B(\MuI._0287_ ),
    .Y(\MuI._0487_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4768_  (.A(\MuI._0286_ ),
    .B(\MuI._0487_ ),
    .Y(\MuI._0488_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4769_  (.A(\MuI._0486_ ),
    .B(\MuI._0488_ ),
    .X(\MuI._0489_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4770_  (.A(\MuI._0465_ ),
    .B(\MuI._0473_ ),
    .C(\MuI._0475_ ),
    .Y(\MuI._0490_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._4771_  (.A1(\MuI._0485_ ),
    .A2(\MuI._0489_ ),
    .B1(\MuI._0490_ ),
    .C1(\MuI._0476_ ),
    .Y(\MuI._0491_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4772_  (.A1(\MuI._0301_ ),
    .A2(\MuI._0302_ ),
    .B1(\MuI._0324_ ),
    .X(\MuI._0492_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4773_  (.A(\MuI._0325_ ),
    .B(\MuI._0492_ ),
    .X(\MuI._0494_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4774_  (.A(\MuI._0476_ ),
    .B(\MuI._0491_ ),
    .C(\MuI._0494_ ),
    .Y(\MuI._0495_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4775_  (.A1(\MuI._0476_ ),
    .A2(\MuI._0491_ ),
    .B1(\MuI._0494_ ),
    .X(\MuI._0496_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._4776_  (.A1(\MuI._0456_ ),
    .A2(\MuI._0495_ ),
    .B1_N(\MuI._0496_ ),
    .X(\MuI._0497_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._4777_  (.A(\MuI._0312_ ),
    .B(\MuI._0313_ ),
    .C(\MuI._0323_ ),
    .Y(\MuI._0498_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4778_  (.A(\MuI._0312_ ),
    .B(\MuI._0498_ ),
    .Y(\MuI._0499_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4779_  (.A(\MuI._0497_ ),
    .B(\MuI._0499_ ),
    .Y(\MuI._0500_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._4780_  (.A1(\MuI._0312_ ),
    .A2(\MuI._0498_ ),
    .B1(\MuI._0497_ ),
    .X(\MuI._0501_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4781_  (.A1(\MuI._0422_ ),
    .A2(\MuI._0500_ ),
    .B1(\MuI._0501_ ),
    .X(\MuI._0502_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4782_  (.A(\MuI.a_operand[19] ),
    .B(\MuI.a_operand[18] ),
    .C(\MuI.b_operand[1] ),
    .D(\MuI.b_operand[0] ),
    .X(\MuI._0503_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4783_  (.A1(\MuI.a_operand[18] ),
    .A2(\MuI._0017_ ),
    .B1(\MuI._0018_ ),
    .B2(\MuI.a_operand[19] ),
    .Y(\MuI._0505_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4784_  (.A_N(\MuI._0503_ ),
    .B_N(\MuI._0505_ ),
    .C(\MuI._2055_ ),
    .D(\MuI._0378_ ),
    .X(\MuI._0506_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4785_  (.A(\MuI._0503_ ),
    .B(\MuI._0506_ ),
    .Y(\MuI._0507_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4786_  (.A1_N(\MuI._1461_ ),
    .A2_N(\MuI._0378_ ),
    .B1(\MuI._0376_ ),
    .B2(\MuI._0377_ ),
    .X(\MuI._0508_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4787_  (.A(\MuI._0379_ ),
    .B(\MuI._0508_ ),
    .Y(\MuI._0509_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4788_  (.A_N(\MuI._0507_ ),
    .B(\MuI._0509_ ),
    .X(\MuI._0510_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4789_  (.A(\MuI._0507_ ),
    .B(\MuI._0509_ ),
    .Y(\MuI._0511_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4790_  (.A(\MuI._0458_ ),
    .B(\MuI._0461_ ),
    .X(\MuI._0512_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4791_  (.A(\MuI._0462_ ),
    .B(\MuI._0512_ ),
    .Y(\MuI._0513_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4792_  (.A(\MuI._0511_ ),
    .B(\MuI._0513_ ),
    .X(\MuI._0514_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4793_  (.A(\MuI._0386_ ),
    .B(\MuI._0388_ ),
    .X(\MuI._0516_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._4794_  (.A1(\MuI._0510_ ),
    .A2(\MuI._0514_ ),
    .B1(\MuI._0516_ ),
    .Y(\MuI._0517_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4795_  (.A(\MuI._0510_ ),
    .B(\MuI._0514_ ),
    .C(\MuI._0516_ ),
    .X(\MuI._0518_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4796_  (.A(\MuI._0469_ ),
    .B(\MuI._0472_ ),
    .Y(\MuI._0519_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4797_  (.A(\MuI._0517_ ),
    .B(\MuI._0518_ ),
    .C(\MuI._0519_ ),
    .Y(\MuI._0520_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4798_  (.A(\MuI._0395_ ),
    .B(\MuI._0392_ ),
    .C(\MuI._0393_ ),
    .X(\MuI._0521_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4799_  (.A1(\MuI._0395_ ),
    .A2(\MuI._0392_ ),
    .B1(\MuI._0393_ ),
    .Y(\MuI._0522_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._4800_  (.A1(\MuI._0517_ ),
    .A2(\MuI._0520_ ),
    .B1(\MuI._0521_ ),
    .C1(\MuI._0522_ ),
    .Y(\MuI._0523_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4801_  (.A1(\MuI._0517_ ),
    .A2(\MuI._0520_ ),
    .B1(\MuI._0521_ ),
    .C1(\MuI._0522_ ),
    .X(\MuI._0524_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4802_  (.A1(\MuI._0521_ ),
    .A2(\MuI._0522_ ),
    .B1(\MuI._0517_ ),
    .C1(\MuI._0520_ ),
    .Y(\MuI._0525_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4803_  (.A1(\MuI._0476_ ),
    .A2(\MuI._0490_ ),
    .B1(\MuI._0489_ ),
    .C1(\MuI._0485_ ),
    .X(\MuI._0527_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4804_  (.A(\MuI._0491_ ),
    .B(\MuI._0524_ ),
    .C(\MuI._0525_ ),
    .D(\MuI._0527_ ),
    .X(\MuI._0528_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4805_  (.A(\MuI._0523_ ),
    .B(\MuI._0528_ ),
    .Y(\MuI._0529_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4806_  (.A(\MuI._0396_ ),
    .B(\MuI._0397_ ),
    .X(\MuI._0530_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4807_  (.A(\MuI._0530_ ),
    .B(\MuI._0399_ ),
    .Y(\MuI._0531_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4808_  (.A(\MuI._0529_ ),
    .B(\MuI._0531_ ),
    .Y(\MuI._0532_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4809_  (.A(\MuI._0496_ ),
    .B(\MuI._0495_ ),
    .X(\MuI._0533_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4810_  (.A(\MuI._0456_ ),
    .B(\MuI._0533_ ),
    .X(\MuI._0534_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4811_  (.A_N(\MuI._0529_ ),
    .B(\MuI._0531_ ),
    .X(\MuI._0535_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4812_  (.A1(\MuI._0532_ ),
    .A2(\MuI._0534_ ),
    .B1(\MuI._0535_ ),
    .Y(\MuI._0536_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4813_  (.A(\MuI._0403_ ),
    .B(\MuI._0404_ ),
    .X(\MuI._0538_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4814_  (.A(\MuI._0536_ ),
    .B(\MuI._0538_ ),
    .Y(\MuI._0539_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4815_  (.A(\MuI._0422_ ),
    .B(\MuI._0500_ ),
    .X(\MuI._0540_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4816_  (.A(\MuI._0536_ ),
    .B_N(\MuI._0538_ ),
    .X(\MuI._0541_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4817_  (.A1(\MuI._0539_ ),
    .A2(\MuI._0540_ ),
    .B1_N(\MuI._0541_ ),
    .Y(\MuI._0542_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4818_  (.A(\MuI._0409_ ),
    .B(\MuI._0410_ ),
    .Y(\MuI._0543_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4819_  (.A(\MuI._0542_ ),
    .B(\MuI._0543_ ),
    .X(\MuI._0544_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4820_  (.A(\MuI._0542_ ),
    .B(\MuI._0543_ ),
    .Y(\MuI._0545_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4821_  (.A1(\MuI._0502_ ),
    .A2(\MuI._0544_ ),
    .B1(\MuI._0545_ ),
    .Y(\MuI._0546_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4822_  (.A(\MuI._0419_ ),
    .B(\MuI._0546_ ),
    .Y(\MuI._0547_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4823_  (.A(\MuI._0285_ ),
    .B(\MuI._0417_ ),
    .X(\MuI._0549_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4824_  (.A(\MuI._0419_ ),
    .B(\MuI._0546_ ),
    .X(\MuI._0550_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4825_  (.A(\MuI._0549_ ),
    .B(\MuI._0550_ ),
    .X(\MuI._0551_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4826_  (.A(\MuI.a_operand[18] ),
    .B(\MuI.a_operand[17] ),
    .C(\MuI.b_operand[1] ),
    .D(\MuI.b_operand[0] ),
    .X(\MuI._0552_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4827_  (.A(\MuI.a_operand[16] ),
    .B(\MuI.b_operand[2] ),
    .Y(\MuI._0553_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4828_  (.A1(\MuI.a_operand[17] ),
    .A2(\MuI.b_operand[1] ),
    .B1(\MuI._0018_ ),
    .B2(\MuI.a_operand[18] ),
    .Y(\MuI._0554_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4829_  (.A(\MuI._0552_ ),
    .B(\MuI._0553_ ),
    .C(\MuI._0554_ ),
    .X(\MuI._0555_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4830_  (.A_N(\MuI._0552_ ),
    .B(\MuI._0555_ ),
    .X(\MuI._0556_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4831_  (.A1_N(\MuI._2843_ ),
    .A2_N(\MuI._3268_ ),
    .B1(\MuI._0503_ ),
    .B2(\MuI._0505_ ),
    .X(\MuI._0557_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4832_  (.A(\MuI._0506_ ),
    .B(\MuI._0557_ ),
    .Y(\MuI._0558_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4833_  (.A_N(\MuI._0556_ ),
    .B(\MuI._0558_ ),
    .X(\MuI._0560_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4834_  (.A(\MuI._0556_ ),
    .B(\MuI._0558_ ),
    .Y(\MuI._0561_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4835_  (.A(\MuI._2671_ ),
    .B(\MuI._2895_ ),
    .Y(\MuI._0562_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4836_  (.A1(\MuI._2605_ ),
    .A2(\MuI._3306_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._2852_ ),
    .Y(\MuI._0563_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4837_  (.A(\MuI._2852_ ),
    .B(\MuI.a_operand[15] ),
    .C(\MuI._2884_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._0564_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4838_  (.A(\MuI._0563_ ),
    .B(\MuI._0564_ ),
    .X(\MuI._0565_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4839_  (.A(\MuI._0562_ ),
    .B(\MuI._0565_ ),
    .Y(\MuI._0566_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4840_  (.A(\MuI._0562_ ),
    .B(\MuI._0565_ ),
    .X(\MuI._0567_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4841_  (.A(\MuI._0566_ ),
    .B(\MuI._0567_ ),
    .Y(\MuI._0568_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4842_  (.A(\MuI._0561_ ),
    .B(\MuI._0568_ ),
    .X(\MuI._0569_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4843_  (.A(\MuI._0511_ ),
    .B(\MuI._0513_ ),
    .X(\MuI._0571_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._4844_  (.A1(\MuI._0560_ ),
    .A2(\MuI._0569_ ),
    .B1(\MuI._0571_ ),
    .Y(\MuI._0572_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4845_  (.A(\MuI._0560_ ),
    .B(\MuI._0569_ ),
    .C(\MuI._0571_ ),
    .X(\MuI._0573_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4846_  (.A(\MuI.a_operand[13] ),
    .B(\MuI.a_operand[12] ),
    .C(\MuI._2866_ ),
    .D(\MuI._2868_ ),
    .X(\MuI._0574_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4847_  (.A1(\MuI._0327_ ),
    .A2(\MuI._3189_ ),
    .B1(\MuI._3190_ ),
    .B2(\MuI._2429_ ),
    .Y(\MuI._0575_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4848_  (.A_N(\MuI._0574_ ),
    .B_N(\MuI._0575_ ),
    .C(\MuI._2484_ ),
    .D(\MuI.b_operand[8] ),
    .X(\MuI._0576_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4849_  (.A(\MuI._0574_ ),
    .B(\MuI._0576_ ),
    .Y(\MuI._0577_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4850_  (.A1_N(\MuI._2451_ ),
    .A2_N(\MuI._0168_ ),
    .B1(\MuI._0466_ ),
    .B2(\MuI._0467_ ),
    .X(\MuI._0578_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4851_  (.A(\MuI._0468_ ),
    .B(\MuI._0578_ ),
    .Y(\MuI._0579_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4852_  (.A1(\MuI._0564_ ),
    .A2(\MuI._0566_ ),
    .B1(\MuI._0579_ ),
    .Y(\MuI._0580_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4853_  (.A(\MuI._0564_ ),
    .B(\MuI._0566_ ),
    .C(\MuI._0579_ ),
    .X(\MuI._0582_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4854_  (.A(\MuI._0580_ ),
    .B(\MuI._0582_ ),
    .X(\MuI._0583_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4855_  (.A(\MuI._0577_ ),
    .B(\MuI._0583_ ),
    .Y(\MuI._0584_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._4856_  (.A(\MuI._0572_ ),
    .B(\MuI._0573_ ),
    .C(\MuI._0584_ ),
    .Y(\MuI._0585_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4857_  (.A1(\MuI._0517_ ),
    .A2(\MuI._0518_ ),
    .B1(\MuI._0519_ ),
    .Y(\MuI._0586_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4858_  (.A(\MuI._0517_ ),
    .B(\MuI._0518_ ),
    .C(\MuI._0519_ ),
    .X(\MuI._0587_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4859_  (.A1(\MuI._0572_ ),
    .A2(\MuI._0585_ ),
    .B1(\MuI._0586_ ),
    .C1(\MuI._0587_ ),
    .X(\MuI._0588_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._4860_  (.A1(\MuI._0572_ ),
    .A2(\MuI._0585_ ),
    .B1(\MuI._0586_ ),
    .C1(\MuI._0587_ ),
    .Y(\MuI._0589_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._4861_  (.A1(\MuI._0587_ ),
    .A2(\MuI._0586_ ),
    .B1(\MuI._0585_ ),
    .C1(\MuI._0572_ ),
    .X(\MuI._0590_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4862_  (.A(\MuI.b_operand[10] ),
    .B(\MuI._2837_ ),
    .C(\MuI.a_operand[10] ),
    .D(\MuI.a_operand[9] ),
    .X(\MuI._0591_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4863_  (.A1(\MuI._2838_ ),
    .A2(\MuI._2765_ ),
    .B1(\MuI._2785_ ),
    .B2(\MuI._2836_ ),
    .Y(\MuI._0593_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4864_  (.A_N(\MuI._0591_ ),
    .B_N(\MuI._0593_ ),
    .C(\MuI._2841_ ),
    .D(\MuI._2352_ ),
    .X(\MuI._0594_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4865_  (.A(\MuI._0591_ ),
    .B(\MuI._0594_ ),
    .Y(\MuI._0595_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4866_  (.A1_N(\MuI._2841_ ),
    .A2_N(\MuI._3223_ ),
    .B1(\MuI._0478_ ),
    .B2(\MuI._0479_ ),
    .X(\MuI._0596_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4867_  (.A(\MuI._0480_ ),
    .B(\MuI._0596_ ),
    .Y(\MuI._0597_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4868_  (.A_N(\MuI._0595_ ),
    .B(\MuI._0597_ ),
    .X(\MuI._0598_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4869_  (.A(\MuI._0597_ ),
    .B(\MuI._0595_ ),
    .Y(\MuI._0599_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4870_  (.A1_N(\MuI._2583_ ),
    .A2_N(\MuI._2330_ ),
    .B1(\MuI._0423_ ),
    .B2(\MuI._0424_ ),
    .X(\MuI._0600_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4871_  (.A(\MuI._0425_ ),
    .B(\MuI._0600_ ),
    .Y(\MuI._0601_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4872_  (.A(\MuI._0599_ ),
    .B(\MuI._0601_ ),
    .X(\MuI._0602_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4873_  (.A(\MuI._0577_ ),
    .B_N(\MuI._0583_ ),
    .X(\MuI._0604_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4874_  (.A(\MuI._0486_ ),
    .B(\MuI._0488_ ),
    .Y(\MuI._0605_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4875_  (.A(\MuI._0489_ ),
    .B(\MuI._0605_ ),
    .X(\MuI._0606_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4876_  (.A1(\MuI._0580_ ),
    .A2(\MuI._0604_ ),
    .B1(\MuI._0606_ ),
    .X(\MuI._0607_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4877_  (.A(\MuI._0580_ ),
    .B(\MuI._0604_ ),
    .C(\MuI._0606_ ),
    .Y(\MuI._0608_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._4878_  (.A1(\MuI._0598_ ),
    .A2(\MuI._0602_ ),
    .B1(\MuI._0607_ ),
    .C1(\MuI._0608_ ),
    .Y(\MuI._0609_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4879_  (.A1(\MuI._0607_ ),
    .A2(\MuI._0608_ ),
    .B1(\MuI._0598_ ),
    .C1(\MuI._0602_ ),
    .X(\MuI._0610_ ));
 sky130_fd_sc_hd__or4bb_1 \MuI._4880_  (.A(\MuI._0589_ ),
    .B(\MuI._0590_ ),
    .C_N(\MuI._0609_ ),
    .D_N(\MuI._0610_ ),
    .X(\MuI._0611_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4881_  (.A1(\MuI._0524_ ),
    .A2(\MuI._0525_ ),
    .B1(\MuI._0527_ ),
    .B2(\MuI._0491_ ),
    .Y(\MuI._0612_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4882_  (.A1(\MuI._0588_ ),
    .A2(\MuI._0611_ ),
    .B1(\MuI._0612_ ),
    .C1(\MuI._0528_ ),
    .X(\MuI._0613_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4883_  (.A1(\MuI._0528_ ),
    .A2(\MuI._0612_ ),
    .B1(\MuI._0611_ ),
    .C1(\MuI._0588_ ),
    .Y(\MuI._0615_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4884_  (.A(\MuI._2799_ ),
    .B(\MuI._2638_ ),
    .C(\MuI._0088_ ),
    .D(\MuI._2319_ ),
    .X(\MuI._0616_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4885_  (.A1(\MuI._2803_ ),
    .A2(\MuI._2374_ ),
    .B1(\MuI._3363_ ),
    .B2(\MuI._2802_ ),
    .Y(\MuI._0617_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4886_  (.A_N(\MuI._0616_ ),
    .B_N(\MuI._0617_ ),
    .C(\MuI._2796_ ),
    .D(\MuI._0101_ ),
    .X(\MuI._0618_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4887_  (.A(\MuI._0616_ ),
    .B(\MuI._0618_ ),
    .Y(\MuI._0619_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4888_  (.A1_N(\MuI._2473_ ),
    .A2_N(\MuI._3372_ ),
    .B1(\MuI._0430_ ),
    .B2(\MuI._0431_ ),
    .X(\MuI._0620_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4889_  (.A(\MuI._0432_ ),
    .B(\MuI._0619_ ),
    .C(\MuI._0620_ ),
    .X(\MuI._0621_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4890_  (.A(\MuI._1296_ ),
    .B(\MuI._1791_ ),
    .C(\MuI._3245_ ),
    .D(\MuI._0304_ ),
    .X(\MuI._0622_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4891_  (.A1(\MuI._2754_ ),
    .A2(\MuI._0228_ ),
    .B1(\MuI._3371_ ),
    .B2(\MuI._3000_ ),
    .Y(\MuI._0623_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4892_  (.A_N(\MuI._0622_ ),
    .B_N(\MuI._0623_ ),
    .C(\MuI._1263_ ),
    .D(\MuI._0445_ ),
    .X(\MuI._0624_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4893_  (.A(\MuI._0622_ ),
    .B(\MuI._0624_ ),
    .X(\MuI._0626_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4894_  (.A(\MuI._0432_ ),
    .B(\MuI._0620_ ),
    .Y(\MuI._0627_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4895_  (.A(\MuI._0619_ ),
    .B(\MuI._0627_ ),
    .Y(\MuI._0628_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4896_  (.A(\MuI._0626_ ),
    .B(\MuI._0628_ ),
    .Y(\MuI._0629_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4897_  (.A(\MuI._0433_ ),
    .B(\MuI._0435_ ),
    .X(\MuI._0630_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4898_  (.A(\MuI._0436_ ),
    .B(\MuI._0630_ ),
    .Y(\MuI._0631_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4899_  (.A1(\MuI._0621_ ),
    .A2(\MuI._0629_ ),
    .B1(\MuI._0631_ ),
    .X(\MuI._0632_ ));
 sky130_fd_sc_hd__inv_2 \MuI._4900_  (.A(\MuI._0632_ ),
    .Y(\MuI._0633_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4901_  (.A(\MuI._0631_ ),
    .B(\MuI._0621_ ),
    .C(\MuI._0629_ ),
    .Y(\MuI._0634_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4902_  (.A(\MuI._0625_ ),
    .B(\MuI._0420_ ),
    .Y(\MuI._0635_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4903_  (.A_N(\MuI._0447_ ),
    .B(\MuI._0446_ ),
    .X(\MuI._0637_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4904_  (.A(\MuI._2817_ ),
    .B(\MuI._0245_ ),
    .Y(\MuI._0638_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4905_  (.A(\MuI._0637_ ),
    .B(\MuI._0638_ ),
    .Y(\MuI._0639_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4906_  (.A(\MuI._2814_ ),
    .B(\MuI._2813_ ),
    .C(\MuI._0111_ ),
    .D(\MuI._0244_ ),
    .X(\MuI._0640_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4907_  (.A1(\MuI._1153_ ),
    .A2(\MuI._0111_ ),
    .B1(\MuI._0315_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._0641_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4908_  (.A_N(\MuI._0640_ ),
    .B_N(\MuI._0641_ ),
    .C(\MuI._2817_ ),
    .D(\MuI._0320_ ),
    .X(\MuI._0642_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4909_  (.A(\MuI._0640_ ),
    .B(\MuI._0642_ ),
    .Y(\MuI._0643_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._4910_  (.A(\MuI._0639_ ),
    .B(\MuI._0643_ ),
    .Y(\MuI._0644_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4911_  (.A(\MuI._0635_ ),
    .B(\MuI._0644_ ),
    .Y(\MuI._0645_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4912_  (.A(\MuI._0632_ ),
    .B(\MuI._0634_ ),
    .C(\MuI._0645_ ),
    .X(\MuI._0646_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4913_  (.A1(\MuI._0440_ ),
    .A2(\MuI._0441_ ),
    .B1(\MuI._0454_ ),
    .Y(\MuI._0648_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4914_  (.A1(\MuI._0607_ ),
    .A2(\MuI._0609_ ),
    .B1(\MuI._0648_ ),
    .C1(\MuI._0455_ ),
    .X(\MuI._0649_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._4915_  (.A1(\MuI._0455_ ),
    .A2(\MuI._0648_ ),
    .B1(\MuI._0609_ ),
    .C1(\MuI._0607_ ),
    .Y(\MuI._0650_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._4916_  (.A1(\MuI._0633_ ),
    .A2(\MuI._0646_ ),
    .B1(\MuI._0649_ ),
    .C1(\MuI._0650_ ),
    .Y(\MuI._0651_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._4917_  (.A1(\MuI._0649_ ),
    .A2(\MuI._0650_ ),
    .B1(\MuI._0633_ ),
    .C1(\MuI._0646_ ),
    .X(\MuI._0652_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._4918_  (.A(\MuI._0613_ ),
    .B(\MuI._0615_ ),
    .C(\MuI._0651_ ),
    .D(\MuI._0652_ ),
    .Y(\MuI._0653_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4919_  (.A(\MuI._0613_ ),
    .B(\MuI._0653_ ),
    .Y(\MuI._0654_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4920_  (.A(\MuI._0532_ ),
    .B(\MuI._0534_ ),
    .X(\MuI._0655_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4921_  (.A(\MuI._0654_ ),
    .B(\MuI._0655_ ),
    .X(\MuI._0656_ ));
 sky130_fd_sc_hd__o22a_1 \MuI._4922_  (.A1(\MuI._0443_ ),
    .A2(\MuI._0448_ ),
    .B1(\MuI._0450_ ),
    .B2(\MuI._0453_ ),
    .X(\MuI._0657_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4923_  (.A1(\MuI._0649_ ),
    .A2(\MuI._0651_ ),
    .B1(\MuI._0657_ ),
    .Y(\MuI._0659_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4924_  (.A(\MuI._0649_ ),
    .B(\MuI._0651_ ),
    .C(\MuI._0657_ ),
    .X(\MuI._0660_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4925_  (.A(\MuI._0659_ ),
    .B(\MuI._0660_ ),
    .Y(\MuI._0661_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._4926_  (.A(\MuI._0452_ ),
    .B(\MuI._0661_ ),
    .X(\MuI._0662_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4927_  (.A(\MuI._0654_ ),
    .B(\MuI._0655_ ),
    .Y(\MuI._0663_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._4928_  (.A1(\MuI._0656_ ),
    .A2(\MuI._0662_ ),
    .B1_N(\MuI._0663_ ),
    .Y(\MuI._0664_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._4929_  (.A(\MuI._0539_ ),
    .B(\MuI._0540_ ),
    .X(\MuI._0665_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4930_  (.A(\MuI._0664_ ),
    .B_N(\MuI._0665_ ),
    .X(\MuI._0666_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4931_  (.A1(\MuI._0452_ ),
    .A2(\MuI._0661_ ),
    .B1(\MuI._0659_ ),
    .X(\MuI._0667_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4932_  (.A(\MuI._0664_ ),
    .B(\MuI._0665_ ),
    .Y(\MuI._0668_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4933_  (.A(\MuI._0667_ ),
    .B(\MuI._0668_ ),
    .Y(\MuI._0670_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4934_  (.A(\MuI._0502_ ),
    .B(\MuI._0544_ ),
    .Y(\MuI._0671_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4935_  (.A1(\MuI._0666_ ),
    .A2(\MuI._0670_ ),
    .B1(\MuI._0671_ ),
    .Y(\MuI._0672_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4936_  (.A(\MuI._0667_ ),
    .B(\MuI._0668_ ),
    .Y(\MuI._0673_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4937_  (.A(\MuI.a_operand[15] ),
    .B(\MuI.a_operand[14] ),
    .C(\MuI._2884_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._0674_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4938_  (.A(\MuI._2440_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._0675_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4939_  (.A1(\MuI._2660_ ),
    .A2(\MuI._2884_ ),
    .B1(\MuI._3307_ ),
    .B2(\MuI._2605_ ),
    .Y(\MuI._0676_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4940_  (.A(\MuI._0674_ ),
    .B(\MuI._0676_ ),
    .X(\MuI._0677_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4941_  (.A(\MuI._0675_ ),
    .B(\MuI._0677_ ),
    .Y(\MuI._0678_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4942_  (.A1_N(\MuI._2484_ ),
    .A2_N(\MuI._0168_ ),
    .B1(\MuI._0574_ ),
    .B2(\MuI._0575_ ),
    .X(\MuI._0679_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4943_  (.A(\MuI._0576_ ),
    .B(\MuI._0679_ ),
    .Y(\MuI._0681_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._4944_  (.A1(\MuI._0674_ ),
    .A2(\MuI._0678_ ),
    .B1(\MuI._0681_ ),
    .Y(\MuI._0682_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4945_  (.A(\MuI.a_operand[12] ),
    .B(\MuI.a_operand[11] ),
    .C(\MuI._2866_ ),
    .D(\MuI._2868_ ),
    .X(\MuI._0683_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4946_  (.A1(\MuI._0477_ ),
    .A2(\MuI._3189_ ),
    .B1(\MuI._3190_ ),
    .B2(\MuI._0327_ ),
    .Y(\MuI._0684_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4947_  (.A_N(\MuI._0683_ ),
    .B_N(\MuI._0684_ ),
    .C(\MuI._2790_ ),
    .D(\MuI.b_operand[8] ),
    .X(\MuI._0685_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4948_  (.A(\MuI._0683_ ),
    .B(\MuI._0685_ ),
    .Y(\MuI._0686_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4949_  (.A(\MuI._0674_ ),
    .B(\MuI._0678_ ),
    .C(\MuI._0681_ ),
    .X(\MuI._0687_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4950_  (.A(\MuI._0682_ ),
    .B(\MuI._0687_ ),
    .X(\MuI._0688_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._4951_  (.A(\MuI._0686_ ),
    .B_N(\MuI._0688_ ),
    .X(\MuI._0689_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4952_  (.A(\MuI._0599_ ),
    .B(\MuI._0601_ ),
    .Y(\MuI._0690_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4953_  (.A(\MuI._0602_ ),
    .B(\MuI._0690_ ),
    .X(\MuI._0692_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._4954_  (.A1(\MuI._0682_ ),
    .A2(\MuI._0689_ ),
    .B1(\MuI._0692_ ),
    .X(\MuI._0693_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4955_  (.A(\MuI.b_operand[10] ),
    .B(\MuI._2837_ ),
    .C(\MuI.a_operand[9] ),
    .D(\MuI.a_operand[8] ),
    .X(\MuI._0694_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4956_  (.A1(\MuI._2837_ ),
    .A2(\MuI.a_operand[9] ),
    .B1(\MuI._2341_ ),
    .B2(\MuI._2853_ ),
    .Y(\MuI._0695_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4957_  (.A_N(\MuI._0694_ ),
    .B_N(\MuI._0695_ ),
    .C(\MuI.b_operand[11] ),
    .D(\MuI._0088_ ),
    .X(\MuI._0696_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4958_  (.A(\MuI._0694_ ),
    .B(\MuI._0696_ ),
    .Y(\MuI._0697_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4959_  (.A1_N(\MuI._2841_ ),
    .A2_N(\MuI._2352_ ),
    .B1(\MuI._0591_ ),
    .B2(\MuI._0593_ ),
    .X(\MuI._0698_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4960_  (.A(\MuI._0594_ ),
    .B(\MuI._0698_ ),
    .Y(\MuI._0699_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4961_  (.A_N(\MuI._0697_ ),
    .B(\MuI._0699_ ),
    .X(\MuI._0700_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4962_  (.A(\MuI._0699_ ),
    .B(\MuI._0697_ ),
    .Y(\MuI._0701_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4963_  (.A1_N(\MuI._2583_ ),
    .A2_N(\MuI._2830_ ),
    .B1(\MuI._0616_ ),
    .B2(\MuI._0617_ ),
    .X(\MuI._0703_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4964_  (.A(\MuI._0618_ ),
    .B(\MuI._0703_ ),
    .Y(\MuI._0704_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4965_  (.A(\MuI._0701_ ),
    .B(\MuI._0704_ ),
    .X(\MuI._0705_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._4966_  (.A(\MuI._0682_ ),
    .B(\MuI._0689_ ),
    .C(\MuI._0692_ ),
    .Y(\MuI._0706_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._4967_  (.A1(\MuI._0700_ ),
    .A2(\MuI._0705_ ),
    .B1(\MuI._0693_ ),
    .C1(\MuI._0706_ ),
    .Y(\MuI._0707_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._4968_  (.A1(\MuI._0632_ ),
    .A2(\MuI._0634_ ),
    .B1(\MuI._0645_ ),
    .Y(\MuI._0708_ ));
 sky130_fd_sc_hd__a211o_2 \MuI._4969_  (.A1(\MuI._0693_ ),
    .A2(\MuI._0707_ ),
    .B1(\MuI._0708_ ),
    .C1(\MuI._0646_ ),
    .X(\MuI._0709_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4970_  (.A(\MuI._2693_ ),
    .B(\MuI._2638_ ),
    .C(\MuI._3362_ ),
    .D(\MuI._0100_ ),
    .X(\MuI._0710_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._4971_  (.A1(\MuI._2918_ ),
    .A2(\MuI._2319_ ),
    .B1(\MuI._2829_ ),
    .B2(\MuI._2799_ ),
    .Y(\MuI._0711_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._4972_  (.A_N(\MuI._0710_ ),
    .B_N(\MuI._0711_ ),
    .C(\MuI.b_operand[14] ),
    .D(\MuI._3246_ ),
    .X(\MuI._0712_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4973_  (.A(\MuI._0710_ ),
    .B(\MuI._0712_ ),
    .Y(\MuI._0714_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4974_  (.A1_N(\MuI._1263_ ),
    .A2_N(\MuI._0445_ ),
    .B1(\MuI._0622_ ),
    .B2(\MuI._0623_ ),
    .X(\MuI._0715_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4975_  (.A(\MuI._0624_ ),
    .B(\MuI._0714_ ),
    .C(\MuI._0715_ ),
    .X(\MuI._0716_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._4976_  (.A1(\MuI._1791_ ),
    .A2(\MuI._0304_ ),
    .B1(\MuI._0444_ ),
    .B2(\MuI._1296_ ),
    .X(\MuI._0717_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4977_  (.A(\MuI._1296_ ),
    .B(\MuI._1791_ ),
    .C(\MuI.a_operand[3] ),
    .D(\MuI._0444_ ),
    .X(\MuI._0718_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._4978_  (.A1(\MuI._1274_ ),
    .A2(\MuI._0245_ ),
    .A3(\MuI._0717_ ),
    .B1(\MuI._0718_ ),
    .X(\MuI._0719_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4979_  (.A(\MuI._0624_ ),
    .B(\MuI._0715_ ),
    .Y(\MuI._0720_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4980_  (.A(\MuI._0714_ ),
    .B(\MuI._0720_ ),
    .Y(\MuI._0721_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4981_  (.A(\MuI._0719_ ),
    .B(\MuI._0721_ ),
    .Y(\MuI._0722_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._4982_  (.A(\MuI._0626_ ),
    .B(\MuI._0628_ ),
    .Y(\MuI._0723_ ));
 sky130_fd_sc_hd__a21oi_4 \MuI._4983_  (.A1(\MuI._0716_ ),
    .A2(\MuI._0722_ ),
    .B1(\MuI._0723_ ),
    .Y(\MuI._0725_ ));
 sky130_fd_sc_hd__and3_1 \MuI._4984_  (.A(\MuI._0723_ ),
    .B(\MuI._0716_ ),
    .C(\MuI._0722_ ),
    .X(\MuI._0726_ ));
 sky130_fd_sc_hd__and4_1 \MuI._4985_  (.A(\MuI._0746_ ),
    .B(\MuI._1164_ ),
    .C(\MuI._0245_ ),
    .D(\MuI._0321_ ),
    .X(\MuI._0727_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._4986_  (.A1_N(\MuI._2817_ ),
    .A2_N(\MuI._0320_ ),
    .B1(\MuI._0640_ ),
    .B2(\MuI._0641_ ),
    .X(\MuI._0728_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4987_  (.A(\MuI._0642_ ),
    .B(\MuI._0728_ ),
    .Y(\MuI._0729_ ));
 sky130_fd_sc_hd__and2_1 \MuI._4988_  (.A(\MuI._0727_ ),
    .B(\MuI._0729_ ),
    .X(\MuI._0730_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._4989_  (.A(\MuI._0727_ ),
    .B(\MuI._0729_ ),
    .Y(\MuI._0731_ ));
 sky130_fd_sc_hd__or2_1 \MuI._4990_  (.A(\MuI._0730_ ),
    .B(\MuI._0731_ ),
    .X(\MuI._0732_ ));
 sky130_fd_sc_hd__or3_1 \MuI._4991_  (.A(\MuI._0725_ ),
    .B(\MuI._0726_ ),
    .C(\MuI._0732_ ),
    .X(\MuI._0733_ ));
 sky130_fd_sc_hd__inv_2 \MuI._4992_  (.A(\MuI._0733_ ),
    .Y(\MuI._0734_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._4993_  (.A1(\MuI._0646_ ),
    .A2(\MuI._0708_ ),
    .B1(\MuI._0707_ ),
    .C1(\MuI._0693_ ),
    .Y(\MuI._0736_ ));
 sky130_fd_sc_hd__o211ai_4 \MuI._4994_  (.A1(\MuI._0725_ ),
    .A2(\MuI._0734_ ),
    .B1(\MuI._0709_ ),
    .C1(\MuI._0736_ ),
    .Y(\MuI._0737_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._4995_  (.A_N(\MuI._0643_ ),
    .B(\MuI._0639_ ),
    .X(\MuI._0738_ ));
 sky130_fd_sc_hd__a31oi_4 \MuI._4996_  (.A1(\MuI._0636_ ),
    .A2(\MuI._0421_ ),
    .A3(\MuI._0644_ ),
    .B1(\MuI._0738_ ),
    .Y(\MuI._0739_ ));
 sky130_fd_sc_hd__a21oi_4 \MuI._4997_  (.A1(\MuI._0709_ ),
    .A2(\MuI._0737_ ),
    .B1(\MuI._0739_ ),
    .Y(\MuI._0740_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._4998_  (.A(\MuI._2605_ ),
    .B(\MuI.b_operand[2] ),
    .Y(\MuI._0741_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._4999_  (.A1(\MuI.a_operand[16] ),
    .A2(\MuI._0017_ ),
    .B1(\MuI._3396_ ),
    .B2(\MuI.a_operand[17] ),
    .Y(\MuI._0742_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5000_  (.A(\MuI.a_operand[17] ),
    .B(\MuI.a_operand[16] ),
    .C(\MuI.b_operand[1] ),
    .D(\MuI.b_operand[0] ),
    .X(\MuI._0743_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5001_  (.A1(\MuI._0741_ ),
    .A2(\MuI._0742_ ),
    .B1_N(\MuI._0743_ ),
    .Y(\MuI._0744_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5002_  (.A1(\MuI._0552_ ),
    .A2(\MuI._0554_ ),
    .B1(\MuI._0553_ ),
    .Y(\MuI._0745_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5003_  (.A(\MuI._0555_ ),
    .B(\MuI._0744_ ),
    .C(\MuI._0745_ ),
    .Y(\MuI._0747_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5004_  (.A1(\MuI._0555_ ),
    .A2(\MuI._0745_ ),
    .B1(\MuI._0744_ ),
    .X(\MuI._0748_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5005_  (.A(\MuI._0675_ ),
    .B(\MuI._0677_ ),
    .X(\MuI._0749_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5006_  (.A(\MuI._0747_ ),
    .B(\MuI._0748_ ),
    .C(\MuI._0749_ ),
    .Y(\MuI._0750_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5007_  (.A(\MuI._0747_ ),
    .B(\MuI._0750_ ),
    .Y(\MuI._0751_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5008_  (.A(\MuI._0561_ ),
    .B(\MuI._0568_ ),
    .X(\MuI._0752_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5009_  (.A(\MuI._0751_ ),
    .B(\MuI._0752_ ),
    .Y(\MuI._0753_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5010_  (.A(\MuI._0753_ ),
    .Y(\MuI._0754_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5011_  (.A(\MuI._0751_ ),
    .B(\MuI._0752_ ),
    .Y(\MuI._0755_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5012_  (.A(\MuI._0686_ ),
    .B(\MuI._0688_ ),
    .Y(\MuI._0756_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5013_  (.A_N(\MuI._0755_ ),
    .B(\MuI._0756_ ),
    .X(\MuI._0758_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5014_  (.A1(\MuI._0572_ ),
    .A2(\MuI._0573_ ),
    .B1(\MuI._0584_ ),
    .X(\MuI._0759_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5015_  (.A1(\MuI._0754_ ),
    .A2(\MuI._0758_ ),
    .B1(\MuI._0759_ ),
    .C1(\MuI._0585_ ),
    .X(\MuI._0760_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5016_  (.A1(\MuI._0585_ ),
    .A2(\MuI._0759_ ),
    .B1(\MuI._0758_ ),
    .C1(\MuI._0754_ ),
    .Y(\MuI._0761_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5017_  (.A1(\MuI._0693_ ),
    .A2(\MuI._0706_ ),
    .B1(\MuI._0700_ ),
    .C1(\MuI._0705_ ),
    .X(\MuI._0762_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._5018_  (.A_N(\MuI._0760_ ),
    .B_N(\MuI._0761_ ),
    .C(\MuI._0707_ ),
    .D(\MuI._0762_ ),
    .X(\MuI._0763_ ));
 sky130_fd_sc_hd__a2bb2o_1 \MuI._5019_  (.A1_N(\MuI._0589_ ),
    .A2_N(\MuI._0590_ ),
    .B1(\MuI._0609_ ),
    .B2(\MuI._0610_ ),
    .X(\MuI._0764_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5020_  (.A1(\MuI._0760_ ),
    .A2(\MuI._0763_ ),
    .B1(\MuI._0764_ ),
    .C1(\MuI._0611_ ),
    .X(\MuI._0765_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5021_  (.A1(\MuI._0611_ ),
    .A2(\MuI._0764_ ),
    .B1(\MuI._0763_ ),
    .C1(\MuI._0760_ ),
    .X(\MuI._0766_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5022_  (.A1(\MuI._0709_ ),
    .A2(\MuI._0736_ ),
    .B1(\MuI._0725_ ),
    .C1(\MuI._0734_ ),
    .X(\MuI._0767_ ));
 sky130_fd_sc_hd__and4b_1 \MuI._5023_  (.A_N(\MuI._0765_ ),
    .B(\MuI._0766_ ),
    .C(\MuI._0737_ ),
    .D(\MuI._0767_ ),
    .X(\MuI._0769_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5024_  (.A1(\MuI._0613_ ),
    .A2(\MuI._0615_ ),
    .B1(\MuI._0651_ ),
    .B2(\MuI._0652_ ),
    .X(\MuI._0770_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5025_  (.A1(\MuI._0765_ ),
    .A2(\MuI._0769_ ),
    .B1(\MuI._0770_ ),
    .C1(\MuI._0653_ ),
    .Y(\MuI._0771_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5026_  (.A1(\MuI._0653_ ),
    .A2(\MuI._0770_ ),
    .B1(\MuI._0769_ ),
    .C1(\MuI._0765_ ),
    .X(\MuI._0772_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5027_  (.A(\MuI._0709_ ),
    .B(\MuI._0737_ ),
    .C(\MuI._0739_ ),
    .X(\MuI._0773_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5028_  (.A(\MuI._0740_ ),
    .B(\MuI._0773_ ),
    .Y(\MuI._0774_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5029_  (.A(\MuI._0771_ ),
    .B(\MuI._0772_ ),
    .C(\MuI._0774_ ),
    .Y(\MuI._0775_ ));
 sky130_fd_sc_hd__and2_2 \MuI._5030_  (.A(\MuI._0771_ ),
    .B(\MuI._0775_ ),
    .X(\MuI._0776_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5031_  (.A(\MuI._0656_ ),
    .B(\MuI._0662_ ),
    .Y(\MuI._0777_ ));
 sky130_fd_sc_hd__xor2_4 \MuI._5032_  (.A(\MuI._0776_ ),
    .B(\MuI._0777_ ),
    .X(\MuI._0778_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5033_  (.A(\MuI._0776_ ),
    .B(\MuI._0777_ ),
    .Y(\MuI._0780_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._5034_  (.A1(\MuI._0740_ ),
    .A2(\MuI._0778_ ),
    .B1(\MuI._0780_ ),
    .Y(\MuI._0781_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5035_  (.A(\MuI._0673_ ),
    .B(\MuI._0781_ ),
    .Y(\MuI._0782_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5036_  (.A(\MuI._0671_ ),
    .B(\MuI._0666_ ),
    .C(\MuI._0670_ ),
    .Y(\MuI._0783_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5037_  (.A1(\MuI._0672_ ),
    .A2(\MuI._0782_ ),
    .B1(\MuI._0783_ ),
    .X(\MuI._0784_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5038_  (.A(\MuI._0285_ ),
    .B(\MuI._0417_ ),
    .Y(\MuI._0785_ ));
 sky130_fd_sc_hd__a221o_1 \MuI._5039_  (.A1(\MuI._0418_ ),
    .A2(\MuI._0547_ ),
    .B1(\MuI._0551_ ),
    .B2(\MuI._0784_ ),
    .C1(\MuI._0785_ ),
    .X(\MuI._0786_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5040_  (.A(\MuI._0148_ ),
    .B(\MuI._0281_ ),
    .Y(\MuI._0787_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5041_  (.A(\MuI._0015_ ),
    .B(\MuI._0139_ ),
    .C(\MuI._0144_ ),
    .Y(\MuI._0788_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._5042_  (.A1(\MuI._0146_ ),
    .A2(\MuI._0787_ ),
    .B1(\MuI._3304_ ),
    .C1(\MuI._0013_ ),
    .D1(\MuI._0788_ ),
    .X(\MuI._0789_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5043_  (.A(\MuI._3305_ ),
    .B(\MuI._0012_ ),
    .X(\MuI._0791_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5044_  (.A1(\MuI._3303_ ),
    .A2(\MuI._0791_ ),
    .B1(\MuI._3302_ ),
    .Y(\MuI._0792_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5045_  (.A1(\MuI._0283_ ),
    .A2(\MuI._0786_ ),
    .B1(\MuI._0789_ ),
    .C1(\MuI._0792_ ),
    .Y(\MuI._0793_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5046_  (.A(\MuI._2799_ ),
    .B(\MuI._2918_ ),
    .C(\MuI.a_operand[1] ),
    .D(\MuI.a_operand[0] ),
    .X(\MuI._0794_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5047_  (.A(\MuI._0794_ ),
    .Y(\MuI._0795_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5048_  (.A(\MuI.a_operand[8] ),
    .B(\MuI.a_operand[7] ),
    .C(\MuI._2884_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._0796_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5049_  (.A1(\MuI._0085_ ),
    .A2(\MuI._3306_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._2341_ ),
    .Y(\MuI._0797_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._5050_  (.A_N(\MuI._0796_ ),
    .B_N(\MuI._0797_ ),
    .C(\MuI._2966_ ),
    .D(\MuI._2319_ ),
    .X(\MuI._0798_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5051_  (.A(\MuI._0796_ ),
    .B(\MuI._0798_ ),
    .Y(\MuI._0799_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5052_  (.A(\MuI._0168_ ),
    .B(\MuI._0228_ ),
    .Y(\MuI._0800_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5053_  (.A(\MuI._3189_ ),
    .B(\MuI._3190_ ),
    .C(\MuI.a_operand[6] ),
    .D(\MuI.a_operand[5] ),
    .X(\MuI._0802_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5054_  (.A1(\MuI._2875_ ),
    .A2(\MuI._3362_ ),
    .B1(\MuI._0100_ ),
    .B2(\MuI._2873_ ),
    .Y(\MuI._0803_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5055_  (.A(\MuI._0802_ ),
    .B(\MuI._0803_ ),
    .Y(\MuI._0804_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5056_  (.A(\MuI._0800_ ),
    .B(\MuI._0804_ ),
    .Y(\MuI._0805_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5057_  (.A(\MuI._0799_ ),
    .B_N(\MuI._0805_ ),
    .X(\MuI._0806_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5058_  (.A(\MuI._2874_ ),
    .B(\MuI._2876_ ),
    .C(\MuI._2830_ ),
    .D(\MuI._3247_ ),
    .X(\MuI._0807_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5059_  (.A(\MuI._2873_ ),
    .B(\MuI._3190_ ),
    .C(\MuI.a_operand[5] ),
    .D(\MuI._3245_ ),
    .Y(\MuI._0808_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5060_  (.A1(\MuI._2868_ ),
    .A2(\MuI.a_operand[5] ),
    .B1(\MuI.a_operand[4] ),
    .B2(\MuI._2866_ ),
    .X(\MuI._0809_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5061_  (.A(\MuI._0168_ ),
    .B(\MuI._3371_ ),
    .C(\MuI._0808_ ),
    .D(\MuI._0809_ ),
    .X(\MuI._0810_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5062_  (.A(\MuI._0807_ ),
    .B(\MuI._0810_ ),
    .Y(\MuI._0811_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5063_  (.A(\MuI._0799_ ),
    .B(\MuI._0805_ ),
    .Y(\MuI._0813_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5064_  (.A(\MuI._0811_ ),
    .B_N(\MuI._0813_ ),
    .X(\MuI._0814_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5065_  (.A(\MuI._2841_ ),
    .B(\MuI._0445_ ),
    .Y(\MuI._0815_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5066_  (.A(\MuI._2853_ ),
    .B(\MuI._2854_ ),
    .C(\MuI.a_operand[4] ),
    .D(\MuI.a_operand[3] ),
    .X(\MuI._0816_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5067_  (.A1(\MuI._2838_ ),
    .A2(\MuI._3245_ ),
    .B1(\MuI._0304_ ),
    .B2(\MuI._2836_ ),
    .Y(\MuI._0817_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5068_  (.A(\MuI._0816_ ),
    .B(\MuI._0817_ ),
    .Y(\MuI._0818_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5069_  (.A(\MuI._0815_ ),
    .B(\MuI._0818_ ),
    .Y(\MuI._0819_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5070_  (.A1(\MuI._2838_ ),
    .A2(\MuI._0304_ ),
    .B1(\MuI._0444_ ),
    .B2(\MuI._2836_ ),
    .X(\MuI._0820_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5071_  (.A(\MuI._2853_ ),
    .B(\MuI._2854_ ),
    .C(\MuI.a_operand[3] ),
    .D(\MuI._0444_ ),
    .X(\MuI._0821_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5072_  (.A1(\MuI._2850_ ),
    .A2(\MuI._0315_ ),
    .A3(\MuI._0820_ ),
    .B1(\MuI._0821_ ),
    .X(\MuI._0822_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5073_  (.A(\MuI._0819_ ),
    .B(\MuI._0822_ ),
    .X(\MuI._0824_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5074_  (.A1(\MuI._2919_ ),
    .A2(\MuI._0315_ ),
    .B1(\MuI.a_operand[0] ),
    .B2(\MuI._2800_ ),
    .X(\MuI._0825_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5075_  (.A(\MuI._0795_ ),
    .B(\MuI._0825_ ),
    .X(\MuI._0826_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5076_  (.A(\MuI._0824_ ),
    .B(\MuI._0826_ ),
    .Y(\MuI._0827_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5077_  (.A1(\MuI._0806_ ),
    .A2(\MuI._0814_ ),
    .B1(\MuI._0827_ ),
    .Y(\MuI._0828_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5078_  (.A(\MuI._2836_ ),
    .B(\MuI._2838_ ),
    .C(\MuI._0444_ ),
    .D(\MuI.a_operand[1] ),
    .X(\MuI._0829_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5079_  (.A1(\MuI._2845_ ),
    .A2(\MuI._0110_ ),
    .B1(\MuI._0244_ ),
    .B2(\MuI._2844_ ),
    .Y(\MuI._0830_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._5080_  (.A_N(\MuI._0829_ ),
    .B_N(\MuI._0830_ ),
    .C(\MuI._2850_ ),
    .D(\MuI.a_operand[0] ),
    .X(\MuI._0831_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5081_  (.A(\MuI._0829_ ),
    .B(\MuI._0831_ ),
    .Y(\MuI._0832_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5082_  (.A(\MuI._2850_ ),
    .B(\MuI._0244_ ),
    .Y(\MuI._0833_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5083_  (.A_N(\MuI._0821_ ),
    .B(\MuI._0820_ ),
    .X(\MuI._0835_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5084_  (.A(\MuI._0833_ ),
    .B(\MuI._0835_ ),
    .Y(\MuI._0836_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5085_  (.A(\MuI._0832_ ),
    .B_N(\MuI._0836_ ),
    .X(\MuI._0837_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5086_  (.A(\MuI._2919_ ),
    .B(\MuI._0321_ ),
    .Y(\MuI._0838_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5087_  (.A(\MuI._0836_ ),
    .B(\MuI._0832_ ),
    .Y(\MuI._0839_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5088_  (.A(\MuI._0838_ ),
    .B_N(\MuI._0839_ ),
    .X(\MuI._0840_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5089_  (.A(\MuI._0806_ ),
    .B(\MuI._0814_ ),
    .C(\MuI._0827_ ),
    .X(\MuI._0841_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5090_  (.A1(\MuI._0837_ ),
    .A2(\MuI._0840_ ),
    .B1(\MuI._0828_ ),
    .C1(\MuI._0841_ ),
    .Y(\MuI._0842_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5091_  (.A(\MuI._0828_ ),
    .B(\MuI._0842_ ),
    .Y(\MuI._0843_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5092_  (.A(\MuI._0795_ ),
    .B(\MuI._0843_ ),
    .X(\MuI._0844_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5093_  (.A(\MuI._0795_ ),
    .B(\MuI._0843_ ),
    .Y(\MuI._0846_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5094_  (.A(\MuI._0844_ ),
    .B(\MuI._0846_ ),
    .X(\MuI._0847_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5095_  (.A(\MuI._2765_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._0848_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5096_  (.A(\MuI.a_operand[12] ),
    .B(\MuI.a_operand[11] ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._0849_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5097_  (.A1(\MuI._0477_ ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._3396_ ),
    .B2(\MuI._0327_ ),
    .Y(\MuI._0850_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5098_  (.A(\MuI._0848_ ),
    .B(\MuI._0849_ ),
    .C(\MuI._0850_ ),
    .X(\MuI._0851_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5099_  (.A1(\MuI._0849_ ),
    .A2(\MuI._0850_ ),
    .B1(\MuI._0848_ ),
    .Y(\MuI._0852_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5100_  (.A(\MuI._2785_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._0853_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5101_  (.A1(\MuI._2765_ ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI._0477_ ),
    .Y(\MuI._0854_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5102_  (.A(\MuI.a_operand[11] ),
    .B(\MuI.a_operand[10] ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._0855_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5103_  (.A1(\MuI._0853_ ),
    .A2(\MuI._0854_ ),
    .B1_N(\MuI._0855_ ),
    .Y(\MuI._0857_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5104_  (.A1(\MuI._0851_ ),
    .A2(\MuI._0852_ ),
    .B1(\MuI._0857_ ),
    .X(\MuI._0858_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5105_  (.A(\MuI._2374_ ),
    .B(\MuI._2895_ ),
    .Y(\MuI._0859_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5106_  (.A1(\MuI._3349_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._3185_ ),
    .B2(\MuI._3223_ ),
    .Y(\MuI._0860_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5107_  (.A(\MuI._2785_ ),
    .B(\MuI._2341_ ),
    .C(\MuI._2885_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._0861_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5108_  (.A(\MuI._0860_ ),
    .B(\MuI._0861_ ),
    .Y(\MuI._0862_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5109_  (.A(\MuI._0859_ ),
    .B(\MuI._0862_ ),
    .Y(\MuI._0863_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5110_  (.A(\MuI._0857_ ),
    .B(\MuI._0851_ ),
    .C(\MuI._0852_ ),
    .Y(\MuI._0864_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5111_  (.A1(\MuI._0858_ ),
    .A2(\MuI._0863_ ),
    .B1_N(\MuI._0864_ ),
    .X(\MuI._0865_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5112_  (.A1(\MuI._2785_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._3185_ ),
    .B2(\MuI._2790_ ),
    .Y(\MuI._0866_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5113_  (.A(\MuI._2765_ ),
    .B(\MuI.a_operand[9] ),
    .C(\MuI._3306_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._0868_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5114_  (.A(\MuI._0866_ ),
    .B(\MuI._0868_ ),
    .Y(\MuI._0869_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5115_  (.A(\MuI._2352_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._0870_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5116_  (.A(\MuI._0869_ ),
    .B(\MuI._0870_ ),
    .Y(\MuI._0871_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5117_  (.A1(\MuI._0848_ ),
    .A2(\MuI._0850_ ),
    .B1_N(\MuI._0849_ ),
    .Y(\MuI._0872_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5118_  (.A(\MuI._0477_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._0873_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5119_  (.A(\MuI.a_operand[13] ),
    .B(\MuI.a_operand[12] ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._0874_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5120_  (.A1(\MuI._0327_ ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._3396_ ),
    .B2(\MuI._2429_ ),
    .Y(\MuI._0875_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5121_  (.A(\MuI._0873_ ),
    .B(\MuI._0874_ ),
    .C(\MuI._0875_ ),
    .X(\MuI._0876_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5122_  (.A1(\MuI._0874_ ),
    .A2(\MuI._0875_ ),
    .B1(\MuI._0873_ ),
    .Y(\MuI._0877_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5123_  (.A(\MuI._0872_ ),
    .B(\MuI._0876_ ),
    .C(\MuI._0877_ ),
    .Y(\MuI._0879_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5124_  (.A1(\MuI._0876_ ),
    .A2(\MuI._0877_ ),
    .B1(\MuI._0872_ ),
    .X(\MuI._0880_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5125_  (.A(\MuI._0871_ ),
    .B(\MuI._0879_ ),
    .C(\MuI._0880_ ),
    .Y(\MuI._0881_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5126_  (.A1(\MuI._0879_ ),
    .A2(\MuI._0880_ ),
    .B1(\MuI._0871_ ),
    .X(\MuI._0882_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5127_  (.A(\MuI._0865_ ),
    .B(\MuI._0881_ ),
    .C(\MuI._0882_ ),
    .Y(\MuI._0883_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5128_  (.A1(\MuI._0881_ ),
    .A2(\MuI._0882_ ),
    .B1(\MuI._0865_ ),
    .X(\MuI._0884_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5129_  (.A1(\MuI._0800_ ),
    .A2(\MuI._0803_ ),
    .B1_N(\MuI._0802_ ),
    .X(\MuI._0885_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5130_  (.A1(\MuI._0859_ ),
    .A2(\MuI._0860_ ),
    .B1_N(\MuI._0861_ ),
    .X(\MuI._0886_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5131_  (.A(\MuI._2871_ ),
    .B(\MuI._0101_ ),
    .Y(\MuI._0887_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5132_  (.A(\MuI._2873_ ),
    .B(\MuI._3190_ ),
    .C(\MuI._0085_ ),
    .D(\MuI.a_operand[6] ),
    .X(\MuI._0888_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5133_  (.A1(\MuI._2869_ ),
    .A2(\MuI._0088_ ),
    .B1(\MuI._2319_ ),
    .B2(\MuI._2867_ ),
    .Y(\MuI._0890_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5134_  (.A(\MuI._0888_ ),
    .B(\MuI._0890_ ),
    .Y(\MuI._0891_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5135_  (.A(\MuI._0887_ ),
    .B(\MuI._0891_ ),
    .Y(\MuI._0892_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5136_  (.A(\MuI._0886_ ),
    .B(\MuI._0892_ ),
    .Y(\MuI._0893_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5137_  (.A(\MuI._0885_ ),
    .B(\MuI._0893_ ),
    .Y(\MuI._0894_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5138_  (.A(\MuI._0883_ ),
    .B(\MuI._0884_ ),
    .C(\MuI._0894_ ),
    .Y(\MuI._0895_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5139_  (.A1(\MuI._0866_ ),
    .A2(\MuI._0870_ ),
    .B1_N(\MuI._0868_ ),
    .X(\MuI._0896_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5140_  (.A(\MuI._0168_ ),
    .B(\MuI._2319_ ),
    .Y(\MuI._0897_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5141_  (.A(\MuI._2866_ ),
    .B(\MuI._2868_ ),
    .C(\MuI.a_operand[8] ),
    .D(\MuI.a_operand[7] ),
    .X(\MuI._0898_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5142_  (.A1(\MuI._2875_ ),
    .A2(\MuI._2341_ ),
    .B1(\MuI._0085_ ),
    .B2(\MuI._2873_ ),
    .Y(\MuI._0899_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5143_  (.A(\MuI._0898_ ),
    .B(\MuI._0899_ ),
    .Y(\MuI._0901_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5144_  (.A(\MuI._0897_ ),
    .B(\MuI._0901_ ),
    .Y(\MuI._0902_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5145_  (.A(\MuI._0896_ ),
    .B(\MuI._0902_ ),
    .Y(\MuI._0903_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5146_  (.A1(\MuI._0887_ ),
    .A2(\MuI._0890_ ),
    .B1_N(\MuI._0888_ ),
    .X(\MuI._0904_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5147_  (.A(\MuI._0903_ ),
    .B(\MuI._0904_ ),
    .Y(\MuI._0905_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5148_  (.A1(\MuI._0871_ ),
    .A2(\MuI._0880_ ),
    .B1_N(\MuI._0879_ ),
    .X(\MuI._0906_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5149_  (.A1(\MuI._2765_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._2484_ ),
    .Y(\MuI._0907_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5150_  (.A(\MuI._0477_ ),
    .B(\MuI._2765_ ),
    .C(\MuI._3306_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._0908_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5151_  (.A(\MuI._0907_ ),
    .B(\MuI._0908_ ),
    .Y(\MuI._0909_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5152_  (.A(\MuI._3223_ ),
    .B(\MuI.b_operand[5] ),
    .Y(\MuI._0910_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5153_  (.A(\MuI._0909_ ),
    .B(\MuI._0910_ ),
    .Y(\MuI._0912_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5154_  (.A1(\MuI._0873_ ),
    .A2(\MuI._0875_ ),
    .B1_N(\MuI._0874_ ),
    .Y(\MuI._0913_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5155_  (.A(\MuI._0327_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._0914_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5156_  (.A(\MuI.a_operand[14] ),
    .B(\MuI.a_operand[13] ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._0915_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5157_  (.A1(\MuI._2429_ ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._3396_ ),
    .B2(\MuI._2660_ ),
    .Y(\MuI._0916_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5158_  (.A(\MuI._0914_ ),
    .B(\MuI._0915_ ),
    .C(\MuI._0916_ ),
    .X(\MuI._0917_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5159_  (.A1(\MuI._0915_ ),
    .A2(\MuI._0916_ ),
    .B1(\MuI._0914_ ),
    .Y(\MuI._0918_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5160_  (.A(\MuI._0913_ ),
    .B(\MuI._0917_ ),
    .C(\MuI._0918_ ),
    .Y(\MuI._0919_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5161_  (.A1(\MuI._0917_ ),
    .A2(\MuI._0918_ ),
    .B1(\MuI._0913_ ),
    .X(\MuI._0920_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5162_  (.A(\MuI._0912_ ),
    .B(\MuI._0919_ ),
    .C(\MuI._0920_ ),
    .Y(\MuI._0921_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5163_  (.A1(\MuI._0919_ ),
    .A2(\MuI._0920_ ),
    .B1(\MuI._0912_ ),
    .X(\MuI._0923_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5164_  (.A(\MuI._0906_ ),
    .B(\MuI._0921_ ),
    .C(\MuI._0923_ ),
    .Y(\MuI._0924_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5165_  (.A1(\MuI._0921_ ),
    .A2(\MuI._0923_ ),
    .B1(\MuI._0906_ ),
    .X(\MuI._0925_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5166_  (.A(\MuI._0905_ ),
    .B(\MuI._0924_ ),
    .C(\MuI._0925_ ),
    .X(\MuI._0926_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5167_  (.A1(\MuI._0924_ ),
    .A2(\MuI._0925_ ),
    .B1(\MuI._0905_ ),
    .Y(\MuI._0927_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._5168_  (.A1(\MuI._0883_ ),
    .A2(\MuI._0895_ ),
    .B1(\MuI._0926_ ),
    .C1(\MuI._0927_ ),
    .Y(\MuI._0928_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5169_  (.A1(\MuI._0926_ ),
    .A2(\MuI._0927_ ),
    .B1(\MuI._0883_ ),
    .C1(\MuI._0895_ ),
    .X(\MuI._0929_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5170_  (.A(\MuI._0886_ ),
    .B_N(\MuI._0892_ ),
    .X(\MuI._0930_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5171_  (.A(\MuI._0885_ ),
    .B_N(\MuI._0893_ ),
    .X(\MuI._0931_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5172_  (.A(\MuI._2841_ ),
    .B(\MuI._0305_ ),
    .Y(\MuI._0932_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5173_  (.A(\MuI._2853_ ),
    .B(\MuI._2854_ ),
    .C(\MuI._0100_ ),
    .D(\MuI._3245_ ),
    .X(\MuI._0934_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5174_  (.A1(\MuI._2838_ ),
    .A2(\MuI._0100_ ),
    .B1(\MuI._0228_ ),
    .B2(\MuI._2844_ ),
    .Y(\MuI._0935_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5175_  (.A(\MuI._0934_ ),
    .B(\MuI._0935_ ),
    .Y(\MuI._0936_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5176_  (.A(\MuI._0932_ ),
    .B(\MuI._0936_ ),
    .Y(\MuI._0937_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5177_  (.A1(\MuI._0815_ ),
    .A2(\MuI._0817_ ),
    .B1_N(\MuI._0816_ ),
    .X(\MuI._0938_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5178_  (.A(\MuI._0937_ ),
    .B(\MuI._0938_ ),
    .Y(\MuI._0939_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5179_  (.A(\MuI._2583_ ),
    .B(\MuI._0320_ ),
    .Y(\MuI._0940_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5180_  (.A(\MuI._2799_ ),
    .B(\MuI._2918_ ),
    .C(\MuI._0110_ ),
    .D(\MuI.a_operand[1] ),
    .X(\MuI._0941_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5181_  (.A1(\MuI._2803_ ),
    .A2(\MuI._0110_ ),
    .B1(\MuI._0244_ ),
    .B2(\MuI._2802_ ),
    .X(\MuI._0942_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5182_  (.A_N(\MuI._0941_ ),
    .B(\MuI._0942_ ),
    .X(\MuI._0943_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5183_  (.A(\MuI._0940_ ),
    .B(\MuI._0943_ ),
    .Y(\MuI._0945_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5184_  (.A(\MuI._0939_ ),
    .B(\MuI._0945_ ),
    .Y(\MuI._0946_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5185_  (.A1(\MuI._0930_ ),
    .A2(\MuI._0931_ ),
    .B1(\MuI._0946_ ),
    .X(\MuI._0947_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5186_  (.A(\MuI._0930_ ),
    .B(\MuI._0931_ ),
    .C(\MuI._0946_ ),
    .Y(\MuI._0948_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5187_  (.A1(\MuI._0819_ ),
    .A2(\MuI._0822_ ),
    .B1(\MuI._0824_ ),
    .B2(\MuI._0826_ ),
    .X(\MuI._0949_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5188_  (.A(\MuI._0947_ ),
    .B(\MuI._0948_ ),
    .C(\MuI._0949_ ),
    .Y(\MuI._0950_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5189_  (.A1(\MuI._0947_ ),
    .A2(\MuI._0948_ ),
    .B1(\MuI._0949_ ),
    .X(\MuI._0951_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._5190_  (.A_N(\MuI._0928_ ),
    .B_N(\MuI._0929_ ),
    .C(\MuI._0950_ ),
    .D(\MuI._0951_ ),
    .X(\MuI._0952_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \MuI._5191_  (.A1_N(\MuI._0928_ ),
    .A2_N(\MuI._0929_ ),
    .B1(\MuI._0950_ ),
    .B2(\MuI._0951_ ),
    .Y(\MuI._0953_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5192_  (.A(\MuI._0853_ ),
    .B(\MuI._0855_ ),
    .C(\MuI._0854_ ),
    .X(\MuI._0954_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5193_  (.A1(\MuI._0855_ ),
    .A2(\MuI._0854_ ),
    .B1(\MuI._0853_ ),
    .Y(\MuI._0956_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5194_  (.A(\MuI._3349_ ),
    .B(\MuI._3268_ ),
    .Y(\MuI._0957_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5195_  (.A1(\MuI._2785_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI._2790_ ),
    .Y(\MuI._0958_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5196_  (.A(\MuI._2765_ ),
    .B(\MuI.a_operand[9] ),
    .C(\MuI._3402_ ),
    .D(\MuI._3396_ ),
    .X(\MuI._0959_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5197_  (.A1(\MuI._0957_ ),
    .A2(\MuI._0958_ ),
    .B1_N(\MuI._0959_ ),
    .Y(\MuI._0960_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5198_  (.A1(\MuI._0954_ ),
    .A2(\MuI._0956_ ),
    .B1(\MuI._0960_ ),
    .X(\MuI._0961_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5199_  (.A1_N(\MuI._2895_ ),
    .A2_N(\MuI._3363_ ),
    .B1(\MuI._0796_ ),
    .B2(\MuI._0797_ ),
    .X(\MuI._0962_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5200_  (.A(\MuI._0798_ ),
    .B(\MuI._0962_ ),
    .Y(\MuI._0963_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5201_  (.A(\MuI._0960_ ),
    .B(\MuI._0954_ ),
    .C(\MuI._0956_ ),
    .Y(\MuI._0964_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5202_  (.A1(\MuI._0961_ ),
    .A2(\MuI._0963_ ),
    .B1_N(\MuI._0964_ ),
    .X(\MuI._0965_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5203_  (.A(\MuI._0864_ ),
    .B(\MuI._0858_ ),
    .C(\MuI._0863_ ),
    .Y(\MuI._0967_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5204_  (.A1(\MuI._0864_ ),
    .A2(\MuI._0858_ ),
    .B1(\MuI._0863_ ),
    .X(\MuI._0968_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5205_  (.A(\MuI._0965_ ),
    .B(\MuI._0967_ ),
    .C(\MuI._0968_ ),
    .Y(\MuI._0969_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5206_  (.A1(\MuI._0967_ ),
    .A2(\MuI._0968_ ),
    .B1(\MuI._0965_ ),
    .X(\MuI._0970_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5207_  (.A(\MuI._0811_ ),
    .B(\MuI._0813_ ),
    .Y(\MuI._0971_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5208_  (.A(\MuI._0969_ ),
    .B(\MuI._0970_ ),
    .C(\MuI._0971_ ),
    .Y(\MuI._0972_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5209_  (.A(\MuI._0883_ ),
    .B(\MuI._0884_ ),
    .C(\MuI._0894_ ),
    .X(\MuI._0973_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5210_  (.A1(\MuI._0883_ ),
    .A2(\MuI._0884_ ),
    .B1(\MuI._0894_ ),
    .Y(\MuI._0974_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5211_  (.A1(\MuI._0969_ ),
    .A2(\MuI._0972_ ),
    .B1(\MuI._0973_ ),
    .C1(\MuI._0974_ ),
    .X(\MuI._0975_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5212_  (.A1(\MuI._0973_ ),
    .A2(\MuI._0974_ ),
    .B1(\MuI._0969_ ),
    .C1(\MuI._0972_ ),
    .Y(\MuI._0976_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5213_  (.A(\MuI._0975_ ),
    .B(\MuI._0976_ ),
    .Y(\MuI._0978_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5214_  (.A1(\MuI._0828_ ),
    .A2(\MuI._0841_ ),
    .B1(\MuI._0837_ ),
    .C1(\MuI._0840_ ),
    .X(\MuI._0979_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5215_  (.A(\MuI._0842_ ),
    .B(\MuI._0979_ ),
    .X(\MuI._0980_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5216_  (.A(\MuI._0978_ ),
    .B(\MuI._0980_ ),
    .X(\MuI._0981_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5217_  (.A1(\MuI._0952_ ),
    .A2(\MuI._0953_ ),
    .B1(\MuI._0975_ ),
    .C1(\MuI._0981_ ),
    .Y(\MuI._0982_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5218_  (.A1(\MuI._0975_ ),
    .A2(\MuI._0981_ ),
    .B1(\MuI._0952_ ),
    .C1(\MuI._0953_ ),
    .X(\MuI._0983_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5219_  (.A1(\MuI._0847_ ),
    .A2(\MuI._0982_ ),
    .B1_N(\MuI._0983_ ),
    .X(\MuI._0984_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5220_  (.A1(\MuI._2860_ ),
    .A2(\MuI._0420_ ),
    .A3(\MuI._0942_ ),
    .B1(\MuI._0941_ ),
    .X(\MuI._0985_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5221_  (.A(\MuI._1813_ ),
    .B(\MuI._0420_ ),
    .C(\MuI._0985_ ),
    .X(\MuI._0986_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5222_  (.A1(\MuI._1813_ ),
    .A2(\MuI._0421_ ),
    .B1(\MuI._0985_ ),
    .Y(\MuI._0987_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5223_  (.A(\MuI._0986_ ),
    .B(\MuI._0987_ ),
    .X(\MuI._0989_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5224_  (.A1(\MuI._0947_ ),
    .A2(\MuI._0950_ ),
    .B1(\MuI._0989_ ),
    .Y(\MuI._0990_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5225_  (.A(\MuI._0947_ ),
    .B(\MuI._0950_ ),
    .C(\MuI._0989_ ),
    .X(\MuI._0991_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5226_  (.A(\MuI._0990_ ),
    .B(\MuI._0991_ ),
    .Y(\MuI._0992_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5227_  (.A(\MuI._0896_ ),
    .B_N(\MuI._0902_ ),
    .X(\MuI._0993_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5228_  (.A(\MuI._0904_ ),
    .B_N(\MuI._0903_ ),
    .X(\MuI._0994_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5229_  (.A(\MuI._2841_ ),
    .B(\MuI._0228_ ),
    .Y(\MuI._0995_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5230_  (.A(\MuI.b_operand[10] ),
    .B(\MuI._2837_ ),
    .C(\MuI.a_operand[6] ),
    .D(\MuI.a_operand[5] ),
    .X(\MuI._0996_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5231_  (.A1(\MuI._2837_ ),
    .A2(\MuI.a_operand[6] ),
    .B1(\MuI.a_operand[5] ),
    .B2(\MuI.b_operand[10] ),
    .X(\MuI._0997_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5232_  (.A_N(\MuI._0996_ ),
    .B(\MuI._0997_ ),
    .X(\MuI._0998_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5233_  (.A(\MuI._0995_ ),
    .B(\MuI._0998_ ),
    .Y(\MuI._1000_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5234_  (.A1(\MuI._0932_ ),
    .A2(\MuI._0935_ ),
    .B1_N(\MuI._0934_ ),
    .X(\MuI._1001_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5235_  (.A(\MuI._1000_ ),
    .B(\MuI._1001_ ),
    .Y(\MuI._1002_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5236_  (.A(\MuI._2583_ ),
    .B(\MuI._0315_ ),
    .Y(\MuI._1003_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5237_  (.A(\MuI._2693_ ),
    .B(\MuI._2638_ ),
    .C(\MuI._0304_ ),
    .D(\MuI._0444_ ),
    .X(\MuI._1004_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5238_  (.A1(\MuI._2918_ ),
    .A2(\MuI._0304_ ),
    .B1(\MuI._0110_ ),
    .B2(\MuI._2799_ ),
    .X(\MuI._1005_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5239_  (.A_N(\MuI._1004_ ),
    .B(\MuI._1005_ ),
    .X(\MuI._1006_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5240_  (.A(\MuI._1003_ ),
    .B(\MuI._1006_ ),
    .Y(\MuI._1007_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5241_  (.A(\MuI._1002_ ),
    .B(\MuI._1007_ ),
    .Y(\MuI._1008_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5242_  (.A1(\MuI._0993_ ),
    .A2(\MuI._0994_ ),
    .B1(\MuI._1008_ ),
    .X(\MuI._1009_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5243_  (.A(\MuI._0993_ ),
    .B(\MuI._0994_ ),
    .C(\MuI._1008_ ),
    .Y(\MuI._1011_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5244_  (.A_N(\MuI._0938_ ),
    .B(\MuI._0937_ ),
    .X(\MuI._1012_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5245_  (.A1(\MuI._0939_ ),
    .A2(\MuI._0945_ ),
    .B1(\MuI._1012_ ),
    .X(\MuI._1013_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5246_  (.A1(\MuI._1009_ ),
    .A2(\MuI._1011_ ),
    .B1(\MuI._1013_ ),
    .Y(\MuI._1014_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5247_  (.A(\MuI._1009_ ),
    .B(\MuI._1011_ ),
    .C(\MuI._1013_ ),
    .X(\MuI._1015_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5248_  (.A(\MuI._0905_ ),
    .B(\MuI._0924_ ),
    .C(\MuI._0925_ ),
    .Y(\MuI._1016_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5249_  (.A1(\MuI._0907_ ),
    .A2(\MuI._0910_ ),
    .B1_N(\MuI._0908_ ),
    .Y(\MuI._1017_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5250_  (.A(\MuI.b_operand[8] ),
    .B(\MuI._0088_ ),
    .Y(\MuI._1018_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5251_  (.A(\MuI._2873_ ),
    .B(\MuI._2785_ ),
    .C(\MuI._2875_ ),
    .D(\MuI._3349_ ),
    .Y(\MuI._1019_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5252_  (.A1(\MuI.a_operand[9] ),
    .A2(\MuI._3190_ ),
    .B1(\MuI._2341_ ),
    .B2(\MuI._3189_ ),
    .X(\MuI._1020_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._5253_  (.A_N(\MuI._1018_ ),
    .B(\MuI._1019_ ),
    .C(\MuI._1020_ ),
    .Y(\MuI._1022_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5254_  (.A1(\MuI._1019_ ),
    .A2(\MuI._1020_ ),
    .B1_N(\MuI._1018_ ),
    .X(\MuI._1023_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5255_  (.A(\MuI._1017_ ),
    .B(\MuI._1022_ ),
    .C(\MuI._1023_ ),
    .Y(\MuI._1024_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5256_  (.A1(\MuI._1022_ ),
    .A2(\MuI._1023_ ),
    .B1(\MuI._1017_ ),
    .X(\MuI._1025_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5257_  (.A1(\MuI._2871_ ),
    .A2(\MuI._2330_ ),
    .A3(\MuI._0901_ ),
    .B1(\MuI._0898_ ),
    .X(\MuI._1026_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5258_  (.A(\MuI._1024_ ),
    .B(\MuI._1025_ ),
    .C(\MuI._1026_ ),
    .X(\MuI._1027_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5259_  (.A1(\MuI._1024_ ),
    .A2(\MuI._1025_ ),
    .B1(\MuI._1026_ ),
    .Y(\MuI._1028_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5260_  (.A(\MuI._1027_ ),
    .B(\MuI._1028_ ),
    .Y(\MuI._1029_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5261_  (.A1(\MuI._0912_ ),
    .A2(\MuI._0920_ ),
    .B1_N(\MuI._0919_ ),
    .X(\MuI._1030_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5262_  (.A(\MuI._0327_ ),
    .B(\MuI._0477_ ),
    .C(\MuI._3306_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._1031_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5263_  (.A1(\MuI._2484_ ),
    .A2(\MuI._2885_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._0327_ ),
    .Y(\MuI._1033_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5264_  (.A(\MuI._1031_ ),
    .B(\MuI._1033_ ),
    .Y(\MuI._1034_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5265_  (.A(\MuI._2773_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._1035_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5266_  (.A(\MuI._1034_ ),
    .B(\MuI._1035_ ),
    .Y(\MuI._1036_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5267_  (.A1(\MuI._0914_ ),
    .A2(\MuI._0916_ ),
    .B1_N(\MuI._0915_ ),
    .Y(\MuI._1037_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5268_  (.A(\MuI._2429_ ),
    .B(\MuI.b_operand[2] ),
    .Y(\MuI._1038_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5269_  (.A(\MuI.a_operand[15] ),
    .B(\MuI.a_operand[14] ),
    .C(\MuI._0017_ ),
    .D(\MuI._0018_ ),
    .X(\MuI._1039_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5270_  (.A1(\MuI.a_operand[14] ),
    .A2(\MuI._3402_ ),
    .B1(\MuI._3396_ ),
    .B2(\MuI.a_operand[15] ),
    .Y(\MuI._1040_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5271_  (.A(\MuI._1038_ ),
    .B(\MuI._1039_ ),
    .C(\MuI._1040_ ),
    .X(\MuI._1041_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5272_  (.A1(\MuI._1039_ ),
    .A2(\MuI._1040_ ),
    .B1(\MuI._1038_ ),
    .Y(\MuI._1042_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5273_  (.A(\MuI._1037_ ),
    .B(\MuI._1041_ ),
    .C(\MuI._1042_ ),
    .Y(\MuI._1044_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5274_  (.A1(\MuI._1041_ ),
    .A2(\MuI._1042_ ),
    .B1(\MuI._1037_ ),
    .X(\MuI._1045_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5275_  (.A(\MuI._1036_ ),
    .B(\MuI._1044_ ),
    .C(\MuI._1045_ ),
    .Y(\MuI._1046_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5276_  (.A1(\MuI._1044_ ),
    .A2(\MuI._1045_ ),
    .B1(\MuI._1036_ ),
    .X(\MuI._1047_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5277_  (.A(\MuI._1030_ ),
    .B(\MuI._1046_ ),
    .C(\MuI._1047_ ),
    .Y(\MuI._1048_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5278_  (.A1(\MuI._1046_ ),
    .A2(\MuI._1047_ ),
    .B1(\MuI._1030_ ),
    .X(\MuI._1049_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5279_  (.A(\MuI._1029_ ),
    .B(\MuI._1048_ ),
    .C(\MuI._1049_ ),
    .X(\MuI._1050_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._5280_  (.A1(\MuI._1048_ ),
    .A2(\MuI._1049_ ),
    .B1(\MuI._1029_ ),
    .Y(\MuI._1051_ ));
 sky130_fd_sc_hd__a211oi_4 \MuI._5281_  (.A1(\MuI._0924_ ),
    .A2(\MuI._1016_ ),
    .B1(\MuI._1050_ ),
    .C1(\MuI._1051_ ),
    .Y(\MuI._1052_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5282_  (.A1(\MuI._1050_ ),
    .A2(\MuI._1051_ ),
    .B1(\MuI._0924_ ),
    .C1(\MuI._1016_ ),
    .X(\MuI._1053_ ));
 sky130_fd_sc_hd__or4_1 \MuI._5283_  (.A(\MuI._1014_ ),
    .B(\MuI._1015_ ),
    .C(\MuI._1052_ ),
    .D(\MuI._1053_ ),
    .X(\MuI._1055_ ));
 sky130_fd_sc_hd__o22ai_1 \MuI._5284_  (.A1(\MuI._1014_ ),
    .A2(\MuI._1015_ ),
    .B1(\MuI._1052_ ),
    .B2(\MuI._1053_ ),
    .Y(\MuI._1056_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5285_  (.A1(\MuI._0928_ ),
    .A2(\MuI._0952_ ),
    .B1(\MuI._1055_ ),
    .C1(\MuI._1056_ ),
    .X(\MuI._1057_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5286_  (.A1(\MuI._1055_ ),
    .A2(\MuI._1056_ ),
    .B1(\MuI._0928_ ),
    .C1(\MuI._0952_ ),
    .X(\MuI._1058_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5287_  (.A(\MuI._1057_ ),
    .B_N(\MuI._1058_ ),
    .X(\MuI._1059_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5288_  (.A(\MuI._0992_ ),
    .B(\MuI._1059_ ),
    .Y(\MuI._1060_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5289_  (.A(\MuI._0984_ ),
    .B(\MuI._1060_ ),
    .Y(\MuI._1061_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5290_  (.A(\MuI._0844_ ),
    .B(\MuI._1061_ ),
    .Y(\MuI._1062_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5291_  (.A(\MuI._2975_ ),
    .B(\MuI._2976_ ),
    .C(\MuI._0245_ ),
    .D(\MuI._0321_ ),
    .X(\MuI._1063_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5292_  (.A1_N(\MuI._2851_ ),
    .A2_N(\MuI._0320_ ),
    .B1(\MuI._0829_ ),
    .B2(\MuI._0830_ ),
    .X(\MuI._1064_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5293_  (.A(\MuI._0831_ ),
    .B(\MuI._1064_ ),
    .Y(\MuI._1066_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5294_  (.A(\MuI._1063_ ),
    .B(\MuI._1066_ ),
    .X(\MuI._1067_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5295_  (.A1(\MuI._2885_ ),
    .A2(\MuI._3362_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._0085_ ),
    .X(\MuI._1068_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5296_  (.A(\MuI._0085_ ),
    .B(\MuI._3306_ ),
    .C(\MuI.a_operand[6] ),
    .D(\MuI._3307_ ),
    .X(\MuI._1069_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5297_  (.A1(\MuI._2967_ ),
    .A2(\MuI._2830_ ),
    .A3(\MuI._1068_ ),
    .B1(\MuI._1069_ ),
    .X(\MuI._1070_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5298_  (.A1(\MuI._0168_ ),
    .A2(\MuI._3371_ ),
    .B1(\MuI._0808_ ),
    .B2(\MuI._0809_ ),
    .X(\MuI._1071_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5299_  (.A_N(\MuI._0810_ ),
    .B(\MuI._1071_ ),
    .X(\MuI._1072_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5300_  (.A(\MuI._1070_ ),
    .B(\MuI._1072_ ),
    .X(\MuI._1073_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5301_  (.A(\MuI._1070_ ),
    .B(\MuI._1072_ ),
    .Y(\MuI._1074_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5302_  (.A1(\MuI._3190_ ),
    .A2(\MuI.a_operand[4] ),
    .B1(\MuI._0304_ ),
    .B2(\MuI._3189_ ),
    .X(\MuI._1075_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5303_  (.A(\MuI._3189_ ),
    .B(\MuI._3190_ ),
    .C(\MuI.a_operand[4] ),
    .D(\MuI.a_operand[3] ),
    .X(\MuI._1077_ ));
 sky130_fd_sc_hd__a31oi_2 \MuI._5304_  (.A1(\MuI._2898_ ),
    .A2(\MuI._0112_ ),
    .A3(\MuI._1075_ ),
    .B1(\MuI._1077_ ),
    .Y(\MuI._1078_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5305_  (.A(\MuI._1074_ ),
    .B(\MuI._1078_ ),
    .Y(\MuI._1079_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5306_  (.A(\MuI._0838_ ),
    .B(\MuI._0839_ ),
    .Y(\MuI._1080_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5307_  (.A1(\MuI._1073_ ),
    .A2(\MuI._1079_ ),
    .B1(\MuI._1080_ ),
    .X(\MuI._1081_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5308_  (.A(\MuI._1073_ ),
    .B(\MuI._1079_ ),
    .C(\MuI._1080_ ),
    .Y(\MuI._1082_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5309_  (.A(\MuI._1081_ ),
    .B(\MuI._1082_ ),
    .Y(\MuI._1083_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5310_  (.A1(\MuI._1067_ ),
    .A2(\MuI._1083_ ),
    .B1(\MuI._1081_ ),
    .X(\MuI._1084_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5311_  (.A(\MuI._0964_ ),
    .B(\MuI._0961_ ),
    .C(\MuI._0963_ ),
    .Y(\MuI._1085_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5312_  (.A1(\MuI._0964_ ),
    .A2(\MuI._0961_ ),
    .B1(\MuI._0963_ ),
    .X(\MuI._1086_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5313_  (.A_N(\MuI._1069_ ),
    .B(\MuI._1068_ ),
    .X(\MuI._1088_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5314_  (.A(\MuI._2895_ ),
    .B(\MuI._0101_ ),
    .Y(\MuI._1089_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5315_  (.A(\MuI._1088_ ),
    .B(\MuI._1089_ ),
    .Y(\MuI._1090_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5316_  (.A(\MuI._0959_ ),
    .B(\MuI._0957_ ),
    .C(\MuI._0958_ ),
    .X(\MuI._1091_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5317_  (.A1(\MuI._0959_ ),
    .A2(\MuI._0958_ ),
    .B1(\MuI._0957_ ),
    .Y(\MuI._1092_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5318_  (.A(\MuI._0088_ ),
    .B(\MuI._3268_ ),
    .Y(\MuI._1093_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5319_  (.A1(\MuI._3349_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._3397_ ),
    .B2(\MuI._2785_ ),
    .Y(\MuI._1094_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5320_  (.A(\MuI._2785_ ),
    .B(\MuI._2341_ ),
    .C(\MuI._3262_ ),
    .D(\MuI._0020_ ),
    .X(\MuI._1095_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5321_  (.A1(\MuI._1093_ ),
    .A2(\MuI._1094_ ),
    .B1_N(\MuI._1095_ ),
    .Y(\MuI._1096_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5322_  (.A1(\MuI._1091_ ),
    .A2(\MuI._1092_ ),
    .B1(\MuI._1096_ ),
    .X(\MuI._1097_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5323_  (.A(\MuI._1091_ ),
    .B(\MuI._1092_ ),
    .C(\MuI._1096_ ),
    .Y(\MuI._1099_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5324_  (.A1(\MuI._1090_ ),
    .A2(\MuI._1097_ ),
    .B1_N(\MuI._1099_ ),
    .X(\MuI._1100_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5325_  (.A(\MuI._1085_ ),
    .B(\MuI._1086_ ),
    .C(\MuI._1100_ ),
    .Y(\MuI._1101_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5326_  (.A(\MuI._1074_ ),
    .B(\MuI._1078_ ),
    .X(\MuI._1102_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5327_  (.A1(\MuI._1085_ ),
    .A2(\MuI._1086_ ),
    .B1(\MuI._1100_ ),
    .X(\MuI._1103_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5328_  (.A(\MuI._1101_ ),
    .B(\MuI._1102_ ),
    .C(\MuI._1103_ ),
    .Y(\MuI._1104_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5329_  (.A(\MuI._0969_ ),
    .B(\MuI._0970_ ),
    .C(\MuI._0971_ ),
    .X(\MuI._1105_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5330_  (.A1(\MuI._0969_ ),
    .A2(\MuI._0970_ ),
    .B1(\MuI._0971_ ),
    .Y(\MuI._1106_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5331_  (.A1(\MuI._1101_ ),
    .A2(\MuI._1104_ ),
    .B1(\MuI._1105_ ),
    .C1(\MuI._1106_ ),
    .Y(\MuI._1107_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5332_  (.A(\MuI._1107_ ),
    .Y(\MuI._1108_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5333_  (.A(\MuI._1067_ ),
    .B(\MuI._1083_ ),
    .Y(\MuI._1110_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5334_  (.A1(\MuI._1105_ ),
    .A2(\MuI._1106_ ),
    .B1(\MuI._1101_ ),
    .C1(\MuI._1104_ ),
    .X(\MuI._1111_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5335_  (.A(\MuI._1107_ ),
    .B(\MuI._1111_ ),
    .X(\MuI._1112_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5336_  (.A(\MuI._1110_ ),
    .B(\MuI._1112_ ),
    .X(\MuI._1113_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5337_  (.A(\MuI._0978_ ),
    .B(\MuI._0980_ ),
    .Y(\MuI._1114_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5338_  (.A(\MuI._0978_ ),
    .B(\MuI._0980_ ),
    .X(\MuI._1115_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5339_  (.A1(\MuI._1108_ ),
    .A2(\MuI._1113_ ),
    .B1(\MuI._1114_ ),
    .C1(\MuI._1115_ ),
    .Y(\MuI._1116_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5340_  (.A1(\MuI._1114_ ),
    .A2(\MuI._1115_ ),
    .B1(\MuI._1108_ ),
    .C1(\MuI._1113_ ),
    .Y(\MuI._1117_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5341_  (.A_N(\MuI._1116_ ),
    .B(\MuI._1117_ ),
    .X(\MuI._1118_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5342_  (.A(\MuI._1084_ ),
    .B(\MuI._1118_ ),
    .Y(\MuI._1119_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5343_  (.A(\MuI._1110_ ),
    .B(\MuI._1112_ ),
    .Y(\MuI._1121_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5344_  (.A(\MuI._1099_ ),
    .B(\MuI._1090_ ),
    .C(\MuI._1097_ ),
    .Y(\MuI._1122_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5345_  (.A1(\MuI._1099_ ),
    .A2(\MuI._1097_ ),
    .B1(\MuI._1090_ ),
    .X(\MuI._1123_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5346_  (.A(\MuI._2892_ ),
    .B(\MuI._2319_ ),
    .C(\MuI._3185_ ),
    .D(\MuI._2829_ ),
    .X(\MuI._1124_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5347_  (.A1(\MuI._3363_ ),
    .A2(\MuI._3185_ ),
    .B1(\MuI._0101_ ),
    .B2(\MuI._2892_ ),
    .Y(\MuI._1125_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5348_  (.A(\MuI._1124_ ),
    .B(\MuI._1125_ ),
    .Y(\MuI._1126_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5349_  (.A(\MuI._2895_ ),
    .B(\MuI._3246_ ),
    .Y(\MuI._1127_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5350_  (.A(\MuI._1126_ ),
    .B(\MuI._1127_ ),
    .Y(\MuI._1128_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5351_  (.A(\MuI._1095_ ),
    .B(\MuI._1093_ ),
    .C(\MuI._1094_ ),
    .X(\MuI._1129_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5352_  (.A1(\MuI._1095_ ),
    .A2(\MuI._1094_ ),
    .B1(\MuI._1093_ ),
    .Y(\MuI._1130_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5353_  (.A(\MuI._3362_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._1132_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5354_  (.A1(\MuI._0085_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI._2341_ ),
    .Y(\MuI._1133_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5355_  (.A(\MuI.a_operand[8] ),
    .B(\MuI.a_operand[7] ),
    .C(\MuI._3402_ ),
    .D(\MuI._3396_ ),
    .X(\MuI._1134_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5356_  (.A1(\MuI._1132_ ),
    .A2(\MuI._1133_ ),
    .B1_N(\MuI._1134_ ),
    .Y(\MuI._1135_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5357_  (.A1(\MuI._1129_ ),
    .A2(\MuI._1130_ ),
    .B1(\MuI._1135_ ),
    .X(\MuI._1136_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5358_  (.A(\MuI._1129_ ),
    .B(\MuI._1130_ ),
    .C(\MuI._1135_ ),
    .Y(\MuI._1137_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5359_  (.A1(\MuI._1128_ ),
    .A2(\MuI._1136_ ),
    .B1_N(\MuI._1137_ ),
    .X(\MuI._1138_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5360_  (.A(\MuI._1122_ ),
    .B(\MuI._1123_ ),
    .C(\MuI._1138_ ),
    .Y(\MuI._1139_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5361_  (.A1(\MuI._1125_ ),
    .A2(\MuI._1127_ ),
    .B1_N(\MuI._1124_ ),
    .X(\MuI._1140_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5362_  (.A(\MuI._2871_ ),
    .B(\MuI._0445_ ),
    .Y(\MuI._1141_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5363_  (.A_N(\MuI._1077_ ),
    .B(\MuI._1075_ ),
    .X(\MuI._1143_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5364_  (.A(\MuI._1141_ ),
    .B(\MuI._1143_ ),
    .Y(\MuI._1144_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5365_  (.A(\MuI._1140_ ),
    .B(\MuI._1144_ ),
    .Y(\MuI._1145_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5366_  (.A(\MuI._2871_ ),
    .B(\MuI._0244_ ),
    .Y(\MuI._1146_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5367_  (.A1(\MuI._2869_ ),
    .A2(\MuI._0305_ ),
    .B1(\MuI._0445_ ),
    .B2(\MuI._2867_ ),
    .Y(\MuI._1147_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5368_  (.A(\MuI._2867_ ),
    .B(\MuI._2869_ ),
    .C(\MuI._3371_ ),
    .D(\MuI._0444_ ),
    .X(\MuI._1148_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5369_  (.A1(\MuI._1146_ ),
    .A2(\MuI._1147_ ),
    .B1_N(\MuI._1148_ ),
    .X(\MuI._1149_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5370_  (.A(\MuI._1145_ ),
    .B(\MuI._1149_ ),
    .Y(\MuI._1150_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5371_  (.A1(\MuI._1122_ ),
    .A2(\MuI._1123_ ),
    .B1(\MuI._1138_ ),
    .X(\MuI._1151_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5372_  (.A(\MuI._1139_ ),
    .B(\MuI._1150_ ),
    .C(\MuI._1151_ ),
    .Y(\MuI._1152_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5373_  (.A(\MuI._1101_ ),
    .B(\MuI._1102_ ),
    .C(\MuI._1103_ ),
    .X(\MuI._1154_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5374_  (.A1(\MuI._1101_ ),
    .A2(\MuI._1103_ ),
    .B1(\MuI._1102_ ),
    .Y(\MuI._1155_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5375_  (.A1(\MuI._1139_ ),
    .A2(\MuI._1152_ ),
    .B1(\MuI._1154_ ),
    .C1(\MuI._1155_ ),
    .X(\MuI._1156_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5376_  (.A(\MuI._1156_ ),
    .Y(\MuI._1157_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5377_  (.A(\MuI._1140_ ),
    .B_N(\MuI._1144_ ),
    .X(\MuI._1158_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5378_  (.A(\MuI._1149_ ),
    .B_N(\MuI._1145_ ),
    .X(\MuI._1159_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5379_  (.A(\MuI._1063_ ),
    .B(\MuI._1066_ ),
    .Y(\MuI._1160_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5380_  (.A1(\MuI._1158_ ),
    .A2(\MuI._1159_ ),
    .B1(\MuI._1160_ ),
    .Y(\MuI._1161_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5381_  (.A(\MuI._1158_ ),
    .B(\MuI._1159_ ),
    .C(\MuI._1160_ ),
    .X(\MuI._1162_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5382_  (.A(\MuI._1161_ ),
    .B(\MuI._1162_ ),
    .Y(\MuI._1163_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5383_  (.A1(\MuI._1154_ ),
    .A2(\MuI._1155_ ),
    .B1(\MuI._1139_ ),
    .C1(\MuI._1152_ ),
    .Y(\MuI._1165_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5384_  (.A(\MuI._1156_ ),
    .B(\MuI._1163_ ),
    .C(\MuI._1165_ ),
    .X(\MuI._1166_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5385_  (.A(\MuI._1157_ ),
    .B(\MuI._1166_ ),
    .Y(\MuI._1167_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5386_  (.A(\MuI._1121_ ),
    .B(\MuI._1167_ ),
    .Y(\MuI._1168_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5387_  (.A(\MuI._1158_ ),
    .B(\MuI._1159_ ),
    .Y(\MuI._1169_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._5388_  (.A(\MuI._1160_ ),
    .B(\MuI._1168_ ),
    .C_N(\MuI._1169_ ),
    .X(\MuI._1170_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5389_  (.A1(\MuI._1121_ ),
    .A2(\MuI._1167_ ),
    .B1(\MuI._1170_ ),
    .X(\MuI._1171_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5390_  (.A(\MuI._1119_ ),
    .B(\MuI._1171_ ),
    .X(\MuI._1172_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5391_  (.A(\MuI._0983_ ),
    .B(\MuI._0847_ ),
    .C(\MuI._0982_ ),
    .X(\MuI._1173_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5392_  (.A1(\MuI._0983_ ),
    .A2(\MuI._0982_ ),
    .B1(\MuI._0847_ ),
    .Y(\MuI._1174_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5393_  (.A(\MuI._1173_ ),
    .B(\MuI._1174_ ),
    .Y(\MuI._1176_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5394_  (.A1(\MuI._1084_ ),
    .A2(\MuI._1117_ ),
    .B1(\MuI._1116_ ),
    .X(\MuI._1177_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5395_  (.A(\MuI._1176_ ),
    .B(\MuI._1177_ ),
    .Y(\MuI._1178_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5396_  (.A(\MuI._1176_ ),
    .B(\MuI._1177_ ),
    .Y(\MuI._1179_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5397_  (.A1(\MuI._1172_ ),
    .A2(\MuI._1178_ ),
    .B1(\MuI._1179_ ),
    .X(\MuI._1180_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5398_  (.A(\MuI._1062_ ),
    .B(\MuI._1180_ ),
    .Y(\MuI._1181_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5399_  (.A(\MuI._1181_ ),
    .Y(\MuI._1182_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5400_  (.A(\MuI._1119_ ),
    .B(\MuI._1171_ ),
    .Y(\MuI._1183_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5401_  (.A(\MuI._1137_ ),
    .B(\MuI._1128_ ),
    .C(\MuI._1136_ ),
    .Y(\MuI._1184_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5402_  (.A1(\MuI._1137_ ),
    .A2(\MuI._1136_ ),
    .B1(\MuI._1128_ ),
    .X(\MuI._1185_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5403_  (.A(\MuI._2892_ ),
    .B(\MuI._2881_ ),
    .C(\MuI._0100_ ),
    .D(\MuI._3245_ ),
    .X(\MuI._1187_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5404_  (.A1(\MuI._3185_ ),
    .A2(\MuI._2829_ ),
    .B1(\MuI._3246_ ),
    .B2(\MuI._2892_ ),
    .Y(\MuI._1188_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5405_  (.A(\MuI._1187_ ),
    .B(\MuI._1188_ ),
    .Y(\MuI._1189_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5406_  (.A(\MuI._2895_ ),
    .B(\MuI._3372_ ),
    .Y(\MuI._1190_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5407_  (.A(\MuI._1189_ ),
    .B(\MuI._1190_ ),
    .Y(\MuI._1191_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5408_  (.A(\MuI._1134_ ),
    .B(\MuI._1132_ ),
    .C(\MuI._1133_ ),
    .X(\MuI._1192_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5409_  (.A1(\MuI._1134_ ),
    .A2(\MuI._1133_ ),
    .B1(\MuI._1132_ ),
    .Y(\MuI._1193_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5410_  (.A(\MuI._0100_ ),
    .B(\MuI._3268_ ),
    .Y(\MuI._1194_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5411_  (.A1(\MuI._3362_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI._0085_ ),
    .Y(\MuI._1195_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5412_  (.A(\MuI.a_operand[7] ),
    .B(\MuI.a_operand[6] ),
    .C(\MuI._3402_ ),
    .D(\MuI._3396_ ),
    .X(\MuI._1196_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5413_  (.A1(\MuI._1194_ ),
    .A2(\MuI._1195_ ),
    .B1_N(\MuI._1196_ ),
    .Y(\MuI._1198_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5414_  (.A1(\MuI._1192_ ),
    .A2(\MuI._1193_ ),
    .B1(\MuI._1198_ ),
    .X(\MuI._1199_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5415_  (.A(\MuI._1192_ ),
    .B(\MuI._1193_ ),
    .C(\MuI._1198_ ),
    .Y(\MuI._1200_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5416_  (.A1(\MuI._1191_ ),
    .A2(\MuI._1199_ ),
    .B1_N(\MuI._1200_ ),
    .X(\MuI._1201_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5417_  (.A(\MuI._1184_ ),
    .B(\MuI._1185_ ),
    .C(\MuI._1201_ ),
    .Y(\MuI._1202_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5418_  (.A1(\MuI._1188_ ),
    .A2(\MuI._1190_ ),
    .B1_N(\MuI._1187_ ),
    .X(\MuI._1203_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5419_  (.A(\MuI._1148_ ),
    .B(\MuI._1147_ ),
    .Y(\MuI._1204_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5420_  (.A(\MuI._1146_ ),
    .B(\MuI._1204_ ),
    .Y(\MuI._1205_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5421_  (.A(\MuI._1203_ ),
    .B(\MuI._1205_ ),
    .Y(\MuI._1206_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5422_  (.A(\MuI._2871_ ),
    .B(\MuI.a_operand[0] ),
    .Y(\MuI._1207_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5423_  (.A1(\MuI._2869_ ),
    .A2(\MuI._0444_ ),
    .B1(\MuI.a_operand[1] ),
    .B2(\MuI._2867_ ),
    .Y(\MuI._1209_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5424_  (.A(\MuI._2873_ ),
    .B(\MuI._2875_ ),
    .C(\MuI._0444_ ),
    .D(\MuI.a_operand[1] ),
    .X(\MuI._1210_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5425_  (.A1(\MuI._1207_ ),
    .A2(\MuI._1209_ ),
    .B1_N(\MuI._1210_ ),
    .X(\MuI._1211_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5426_  (.A(\MuI._1206_ ),
    .B(\MuI._1211_ ),
    .Y(\MuI._1212_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5427_  (.A1(\MuI._1184_ ),
    .A2(\MuI._1185_ ),
    .B1(\MuI._1201_ ),
    .X(\MuI._1213_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5428_  (.A(\MuI._1202_ ),
    .B(\MuI._1212_ ),
    .C(\MuI._1213_ ),
    .Y(\MuI._1214_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5429_  (.A(\MuI._1139_ ),
    .B(\MuI._1150_ ),
    .C(\MuI._1151_ ),
    .X(\MuI._1215_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5430_  (.A1(\MuI._1139_ ),
    .A2(\MuI._1151_ ),
    .B1(\MuI._1150_ ),
    .Y(\MuI._1216_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5431_  (.A1(\MuI._1202_ ),
    .A2(\MuI._1214_ ),
    .B1(\MuI._1215_ ),
    .C1(\MuI._1216_ ),
    .X(\MuI._1217_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5432_  (.A(\MuI._1203_ ),
    .B_N(\MuI._1205_ ),
    .X(\MuI._1218_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5433_  (.A(\MuI._1211_ ),
    .B_N(\MuI._1206_ ),
    .X(\MuI._1220_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5434_  (.A1(\MuI._2976_ ),
    .A2(\MuI._0246_ ),
    .B1(\MuI._0321_ ),
    .B2(\MuI._2975_ ),
    .Y(\MuI._1221_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5435_  (.A(\MuI._1063_ ),
    .B(\MuI._1221_ ),
    .X(\MuI._1222_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5436_  (.A1(\MuI._1218_ ),
    .A2(\MuI._1220_ ),
    .B1(\MuI._1222_ ),
    .Y(\MuI._1223_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5437_  (.A(\MuI._1218_ ),
    .B(\MuI._1220_ ),
    .C(\MuI._1222_ ),
    .X(\MuI._1224_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5438_  (.A(\MuI._1223_ ),
    .B(\MuI._1224_ ),
    .Y(\MuI._1225_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5439_  (.A1(\MuI._1215_ ),
    .A2(\MuI._1216_ ),
    .B1(\MuI._1202_ ),
    .C1(\MuI._1214_ ),
    .Y(\MuI._1226_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5440_  (.A(\MuI._1217_ ),
    .B(\MuI._1225_ ),
    .C(\MuI._1226_ ),
    .Y(\MuI._1227_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5441_  (.A1(\MuI._1156_ ),
    .A2(\MuI._1165_ ),
    .B1(\MuI._1163_ ),
    .Y(\MuI._1228_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._5442_  (.A1(\MuI._1217_ ),
    .A2(\MuI._1227_ ),
    .B1(\MuI._1166_ ),
    .C1(\MuI._1228_ ),
    .Y(\MuI._1229_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5443_  (.A1(\MuI._1217_ ),
    .A2(\MuI._1227_ ),
    .B1(\MuI._1166_ ),
    .C1(\MuI._1228_ ),
    .X(\MuI._1231_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5444_  (.A1(\MuI._1166_ ),
    .A2(\MuI._1228_ ),
    .B1(\MuI._1217_ ),
    .C1(\MuI._1227_ ),
    .Y(\MuI._1232_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5445_  (.A(\MuI._1223_ ),
    .B(\MuI._1231_ ),
    .C(\MuI._1232_ ),
    .X(\MuI._1233_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5446_  (.A(\MuI._1161_ ),
    .B(\MuI._1168_ ),
    .Y(\MuI._1234_ ));
 sky130_fd_sc_hd__o21ai_4 \MuI._5447_  (.A1(\MuI._1229_ ),
    .A2(\MuI._1233_ ),
    .B1(\MuI._1234_ ),
    .Y(\MuI._1235_ ));
 sky130_fd_sc_hd__nor3_2 \MuI._5448_  (.A(\MuI._1178_ ),
    .B(\MuI._1183_ ),
    .C(\MuI._1235_ ),
    .Y(\MuI._1236_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5449_  (.A1(\MuI._1183_ ),
    .A2(\MuI._1235_ ),
    .B1(\MuI._1172_ ),
    .X(\MuI._1237_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5450_  (.A(\MuI._1178_ ),
    .B(\MuI._1237_ ),
    .Y(\MuI._1238_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5451_  (.A(\MuI._1181_ ),
    .B(\MuI._1238_ ),
    .Y(\MuI._1239_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5452_  (.A(\MuI._1234_ ),
    .B(\MuI._1229_ ),
    .C(\MuI._1233_ ),
    .X(\MuI._1240_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5453_  (.A(\MuI._1235_ ),
    .B(\MuI._1240_ ),
    .Y(\MuI._1242_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5454_  (.A(\MuI._1200_ ),
    .B(\MuI._1191_ ),
    .C(\MuI._1199_ ),
    .Y(\MuI._1243_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5455_  (.A1(\MuI._1200_ ),
    .A2(\MuI._1199_ ),
    .B1(\MuI._1191_ ),
    .X(\MuI._1244_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5456_  (.A1(\MuI._2881_ ),
    .A2(\MuI._3245_ ),
    .B1(\MuI._0304_ ),
    .B2(\MuI._2892_ ),
    .Y(\MuI._1245_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5457_  (.A(\MuI._3306_ ),
    .B(\MuI._3307_ ),
    .C(\MuI.a_operand[4] ),
    .D(\MuI.a_operand[3] ),
    .X(\MuI._1246_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5458_  (.A(\MuI._1245_ ),
    .B(\MuI._1246_ ),
    .Y(\MuI._1247_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5459_  (.A(\MuI._2895_ ),
    .B(\MuI._0111_ ),
    .Y(\MuI._1248_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5460_  (.A(\MuI._1247_ ),
    .B(\MuI._1248_ ),
    .Y(\MuI._1249_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5461_  (.A(\MuI._1196_ ),
    .B(\MuI._1194_ ),
    .C(\MuI._1195_ ),
    .X(\MuI._1250_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5462_  (.A1(\MuI._1196_ ),
    .A2(\MuI._1195_ ),
    .B1(\MuI._1194_ ),
    .Y(\MuI._1251_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5463_  (.A(\MuI._3268_ ),
    .B(\MuI._0228_ ),
    .Y(\MuI._1253_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5464_  (.A1(\MuI._0100_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._3397_ ),
    .B2(\MuI._3362_ ),
    .Y(\MuI._1254_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5465_  (.A(\MuI.a_operand[6] ),
    .B(\MuI.a_operand[5] ),
    .C(\MuI._3262_ ),
    .D(\MuI._0020_ ),
    .X(\MuI._1255_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5466_  (.A1(\MuI._1253_ ),
    .A2(\MuI._1254_ ),
    .B1_N(\MuI._1255_ ),
    .Y(\MuI._1256_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5467_  (.A1(\MuI._1250_ ),
    .A2(\MuI._1251_ ),
    .B1(\MuI._1256_ ),
    .X(\MuI._1257_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5468_  (.A(\MuI._1250_ ),
    .B(\MuI._1251_ ),
    .C(\MuI._1256_ ),
    .Y(\MuI._1258_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5469_  (.A1(\MuI._1249_ ),
    .A2(\MuI._1257_ ),
    .B1_N(\MuI._1258_ ),
    .X(\MuI._1259_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5470_  (.A(\MuI._1243_ ),
    .B(\MuI._1244_ ),
    .C(\MuI._1259_ ),
    .Y(\MuI._1260_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5471_  (.A1(\MuI._2967_ ),
    .A2(\MuI._0111_ ),
    .A3(\MuI._1247_ ),
    .B1(\MuI._1246_ ),
    .X(\MuI._1261_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5472_  (.A(\MuI._1210_ ),
    .B(\MuI._1209_ ),
    .Y(\MuI._1262_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5473_  (.A(\MuI._1207_ ),
    .B(\MuI._1262_ ),
    .Y(\MuI._1264_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5474_  (.A(\MuI._1261_ ),
    .B(\MuI._1264_ ),
    .X(\MuI._1265_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5475_  (.A(\MuI._2874_ ),
    .B(\MuI._2876_ ),
    .C(\MuI._0315_ ),
    .D(\MuI.a_operand[0] ),
    .X(\MuI._1266_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5476_  (.A(\MuI._1265_ ),
    .B(\MuI._1266_ ),
    .X(\MuI._1267_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5477_  (.A1(\MuI._1243_ ),
    .A2(\MuI._1244_ ),
    .B1(\MuI._1259_ ),
    .X(\MuI._1268_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5478_  (.A(\MuI._1260_ ),
    .B(\MuI._1267_ ),
    .C(\MuI._1268_ ),
    .Y(\MuI._1269_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5479_  (.A(\MuI._1202_ ),
    .B(\MuI._1212_ ),
    .C(\MuI._1213_ ),
    .X(\MuI._1270_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._5480_  (.A1(\MuI._1202_ ),
    .A2(\MuI._1213_ ),
    .B1(\MuI._1212_ ),
    .Y(\MuI._1271_ ));
 sky130_fd_sc_hd__a211oi_4 \MuI._5481_  (.A1(\MuI._1260_ ),
    .A2(\MuI._1269_ ),
    .B1(\MuI._1270_ ),
    .C1(\MuI._1271_ ),
    .Y(\MuI._1272_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5482_  (.A(\MuI._1261_ ),
    .B(\MuI._1264_ ),
    .X(\MuI._1273_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5483_  (.A(\MuI._1265_ ),
    .B(\MuI._1266_ ),
    .X(\MuI._1275_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5484_  (.A1(\MuI._1273_ ),
    .A2(\MuI._1275_ ),
    .B1(\MuI._2976_ ),
    .C1(\MuI._0420_ ),
    .X(\MuI._1276_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5485_  (.A1(\MuI._2976_ ),
    .A2(\MuI._0421_ ),
    .B1(\MuI._1273_ ),
    .C1(\MuI._1275_ ),
    .Y(\MuI._1277_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5486_  (.A(\MuI._1276_ ),
    .B(\MuI._1277_ ),
    .X(\MuI._1278_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5487_  (.A1(\MuI._1270_ ),
    .A2(\MuI._1271_ ),
    .B1(\MuI._1260_ ),
    .C1(\MuI._1269_ ),
    .X(\MuI._1279_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5488_  (.A(\MuI._1272_ ),
    .B(\MuI._1278_ ),
    .C(\MuI._1279_ ),
    .Y(\MuI._1280_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5489_  (.A1(\MuI._1217_ ),
    .A2(\MuI._1226_ ),
    .B1(\MuI._1225_ ),
    .X(\MuI._1281_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5490_  (.A1(\MuI._1272_ ),
    .A2(\MuI._1280_ ),
    .B1(\MuI._1227_ ),
    .C1(\MuI._1281_ ),
    .Y(\MuI._1282_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5491_  (.A1(\MuI._1227_ ),
    .A2(\MuI._1281_ ),
    .B1(\MuI._1272_ ),
    .C1(\MuI._1280_ ),
    .X(\MuI._1283_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5492_  (.A(\MuI._1276_ ),
    .B(\MuI._1282_ ),
    .C(\MuI._1283_ ),
    .Y(\MuI._1284_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5493_  (.A1(\MuI._1231_ ),
    .A2(\MuI._1232_ ),
    .B1(\MuI._1223_ ),
    .Y(\MuI._1286_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5494_  (.A1(\MuI._1282_ ),
    .A2(\MuI._1284_ ),
    .B1(\MuI._1233_ ),
    .C1(\MuI._1286_ ),
    .X(\MuI._1287_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5495_  (.A(\MuI._1183_ ),
    .B(\MuI._1242_ ),
    .C(\MuI._1287_ ),
    .X(\MuI._1288_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5496_  (.A1(\MuI._1242_ ),
    .A2(\MuI._1287_ ),
    .B1(\MuI._1183_ ),
    .C1(\MuI._1235_ ),
    .Y(\MuI._1289_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5497_  (.A1(\MuI._1183_ ),
    .A2(\MuI._1235_ ),
    .B1(\MuI._1288_ ),
    .C1(\MuI._1289_ ),
    .Y(\MuI._1290_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5498_  (.A1(\MuI._1233_ ),
    .A2(\MuI._1286_ ),
    .B1(\MuI._1282_ ),
    .C1(\MuI._1284_ ),
    .Y(\MuI._1291_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5499_  (.A(\MuI._1276_ ),
    .B(\MuI._1282_ ),
    .C(\MuI._1283_ ),
    .X(\MuI._1292_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5500_  (.A1(\MuI._1282_ ),
    .A2(\MuI._1283_ ),
    .B1(\MuI._1276_ ),
    .Y(\MuI._1293_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5501_  (.A(\MuI._1292_ ),
    .B(\MuI._1293_ ),
    .Y(\MuI._1294_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5502_  (.A(\MuI._1258_ ),
    .B(\MuI._1249_ ),
    .C(\MuI._1257_ ),
    .Y(\MuI._1295_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5503_  (.A1(\MuI._1258_ ),
    .A2(\MuI._1257_ ),
    .B1(\MuI._1249_ ),
    .X(\MuI._1297_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5504_  (.A1(\MuI._2882_ ),
    .A2(\MuI._0305_ ),
    .B1(\MuI._0445_ ),
    .B2(\MuI._2886_ ),
    .Y(\MuI._1298_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5505_  (.A(\MuI._2892_ ),
    .B(\MuI._3185_ ),
    .C(\MuI._3371_ ),
    .D(\MuI._0110_ ),
    .X(\MuI._1299_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5506_  (.A(\MuI._1298_ ),
    .B(\MuI._1299_ ),
    .Y(\MuI._1300_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5507_  (.A(\MuI._2967_ ),
    .B(\MuI._0315_ ),
    .Y(\MuI._1301_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5508_  (.A(\MuI._1300_ ),
    .B(\MuI._1301_ ),
    .Y(\MuI._1302_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5509_  (.A(\MuI._1255_ ),
    .B(\MuI._1253_ ),
    .C(\MuI._1254_ ),
    .X(\MuI._1303_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5510_  (.A1(\MuI._1255_ ),
    .A2(\MuI._1254_ ),
    .B1(\MuI._1253_ ),
    .Y(\MuI._1304_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5511_  (.A(\MuI._3268_ ),
    .B(\MuI._3371_ ),
    .Y(\MuI._1305_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5512_  (.A1(\MuI._3403_ ),
    .A2(\MuI._3245_ ),
    .B1(\MuI._3397_ ),
    .B2(\MuI._0100_ ),
    .Y(\MuI._1306_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5513_  (.A(\MuI._0100_ ),
    .B(\MuI._3262_ ),
    .C(\MuI.a_operand[4] ),
    .D(\MuI._0020_ ),
    .X(\MuI._1308_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5514_  (.A1(\MuI._1305_ ),
    .A2(\MuI._1306_ ),
    .B1_N(\MuI._1308_ ),
    .Y(\MuI._1309_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5515_  (.A1(\MuI._1303_ ),
    .A2(\MuI._1304_ ),
    .B1(\MuI._1309_ ),
    .X(\MuI._1310_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5516_  (.A(\MuI._1303_ ),
    .B(\MuI._1304_ ),
    .C(\MuI._1309_ ),
    .Y(\MuI._1311_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5517_  (.A1(\MuI._1302_ ),
    .A2(\MuI._1310_ ),
    .B1_N(\MuI._1311_ ),
    .X(\MuI._1312_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5518_  (.A(\MuI._1295_ ),
    .B(\MuI._1297_ ),
    .C(\MuI._1312_ ),
    .Y(\MuI._1313_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5519_  (.A1(\MuI._2967_ ),
    .A2(\MuI._0245_ ),
    .A3(\MuI._1300_ ),
    .B1(\MuI._1299_ ),
    .X(\MuI._1314_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5520_  (.A1(\MuI._2876_ ),
    .A2(\MuI._0245_ ),
    .B1(\MuI._0320_ ),
    .B2(\MuI._2874_ ),
    .Y(\MuI._1315_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5521_  (.A(\MuI._1266_ ),
    .B(\MuI._1315_ ),
    .X(\MuI._1316_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5522_  (.A(\MuI._1314_ ),
    .B(\MuI._1316_ ),
    .Y(\MuI._1317_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5523_  (.A1(\MuI._1295_ ),
    .A2(\MuI._1297_ ),
    .B1(\MuI._1312_ ),
    .X(\MuI._1319_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5524_  (.A(\MuI._1313_ ),
    .B(\MuI._1317_ ),
    .C(\MuI._1319_ ),
    .Y(\MuI._1320_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5525_  (.A(\MuI._1260_ ),
    .B(\MuI._1267_ ),
    .C(\MuI._1268_ ),
    .X(\MuI._1321_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5526_  (.A1(\MuI._1260_ ),
    .A2(\MuI._1268_ ),
    .B1(\MuI._1267_ ),
    .Y(\MuI._1322_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._5527_  (.A1(\MuI._1313_ ),
    .A2(\MuI._1320_ ),
    .B1(\MuI._1321_ ),
    .C1(\MuI._1322_ ),
    .Y(\MuI._1323_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5528_  (.A1(\MuI._1321_ ),
    .A2(\MuI._1322_ ),
    .B1(\MuI._1313_ ),
    .C1(\MuI._1320_ ),
    .X(\MuI._1324_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5529_  (.A_N(\MuI._1316_ ),
    .B(\MuI._1314_ ),
    .X(\MuI._1325_ ));
 sky130_fd_sc_hd__nor3b_1 \MuI._5530_  (.A(\MuI._1323_ ),
    .B(\MuI._1324_ ),
    .C_N(\MuI._1325_ ),
    .Y(\MuI._1326_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5531_  (.A(\MuI._1272_ ),
    .B(\MuI._1278_ ),
    .C(\MuI._1279_ ),
    .X(\MuI._1327_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5532_  (.A1(\MuI._1272_ ),
    .A2(\MuI._1279_ ),
    .B1(\MuI._1278_ ),
    .Y(\MuI._1328_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5533_  (.A1(\MuI._1323_ ),
    .A2(\MuI._1326_ ),
    .B1(\MuI._1327_ ),
    .C1(\MuI._1328_ ),
    .X(\MuI._1330_ ));
 sky130_fd_sc_hd__nand4_2 \MuI._5534_  (.A(\MuI._1287_ ),
    .B(\MuI._1291_ ),
    .C(\MuI._1294_ ),
    .D(\MuI._1330_ ),
    .Y(\MuI._1331_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5535_  (.A1(\MuI._1287_ ),
    .A2(\MuI._1291_ ),
    .B1(\MuI._1294_ ),
    .B2(\MuI._1330_ ),
    .X(\MuI._1332_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5536_  (.A1(\MuI._1327_ ),
    .A2(\MuI._1328_ ),
    .B1(\MuI._1323_ ),
    .C1(\MuI._1326_ ),
    .X(\MuI._1333_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5537_  (.A(\MuI._1330_ ),
    .B_N(\MuI._1333_ ),
    .X(\MuI._1334_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5538_  (.A(\MuI._2886_ ),
    .B(\MuI._2882_ ),
    .C(\MuI._0111_ ),
    .D(\MuI._0315_ ),
    .X(\MuI._1335_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5539_  (.A1(\MuI._3185_ ),
    .A2(\MuI._0110_ ),
    .B1(\MuI.a_operand[1] ),
    .B2(\MuI._2892_ ),
    .X(\MuI._1336_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5540_  (.A(\MuI._2886_ ),
    .B(\MuI._2882_ ),
    .C(\MuI._0445_ ),
    .D(\MuI._0244_ ),
    .Y(\MuI._1337_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5541_  (.A(\MuI._2966_ ),
    .B(\MuI.a_operand[0] ),
    .X(\MuI._1338_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5542_  (.A(\MuI._1336_ ),
    .B(\MuI._1337_ ),
    .C(\MuI._1338_ ),
    .X(\MuI._1339_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5543_  (.A1(\MuI._1335_ ),
    .A2(\MuI._1339_ ),
    .B1(\MuI._2876_ ),
    .C1(\MuI._0321_ ),
    .X(\MuI._1341_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5544_  (.A1(\MuI._2876_ ),
    .A2(\MuI._0321_ ),
    .B1(\MuI._1335_ ),
    .C1(\MuI._1339_ ),
    .Y(\MuI._1342_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5545_  (.A(\MuI._1341_ ),
    .B(\MuI._1342_ ),
    .X(\MuI._1343_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5546_  (.A(\MuI._1311_ ),
    .B(\MuI._1302_ ),
    .C(\MuI._1310_ ),
    .Y(\MuI._1344_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5547_  (.A1(\MuI._1311_ ),
    .A2(\MuI._1310_ ),
    .B1(\MuI._1302_ ),
    .X(\MuI._1345_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5548_  (.A1(\MuI._1336_ ),
    .A2(\MuI._1337_ ),
    .B1(\MuI._1338_ ),
    .Y(\MuI._1346_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5549_  (.A(\MuI._1346_ ),
    .B(\MuI._1339_ ),
    .Y(\MuI._1347_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5550_  (.A(\MuI._1308_ ),
    .B(\MuI._1305_ ),
    .C(\MuI._1306_ ),
    .X(\MuI._1348_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5551_  (.A1(\MuI._1308_ ),
    .A2(\MuI._1306_ ),
    .B1(\MuI._1305_ ),
    .Y(\MuI._1349_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5552_  (.A(\MuI._3268_ ),
    .B(\MuI._0445_ ),
    .Y(\MuI._1350_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5553_  (.A1(\MuI._0228_ ),
    .A2(\MuI._3397_ ),
    .B1(\MuI._0305_ ),
    .B2(\MuI._3403_ ),
    .Y(\MuI._1352_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5554_  (.A(\MuI._3403_ ),
    .B(\MuI._3245_ ),
    .C(\MuI._0020_ ),
    .D(\MuI._0304_ ),
    .X(\MuI._1353_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5555_  (.A1(\MuI._1350_ ),
    .A2(\MuI._1352_ ),
    .B1_N(\MuI._1353_ ),
    .Y(\MuI._1354_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5556_  (.A1(\MuI._1348_ ),
    .A2(\MuI._1349_ ),
    .B1(\MuI._1354_ ),
    .X(\MuI._1355_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5557_  (.A(\MuI._1348_ ),
    .B(\MuI._1349_ ),
    .C(\MuI._1354_ ),
    .Y(\MuI._1356_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5558_  (.A1(\MuI._1347_ ),
    .A2(\MuI._1355_ ),
    .B1_N(\MuI._1356_ ),
    .X(\MuI._1357_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5559_  (.A1(\MuI._1344_ ),
    .A2(\MuI._1345_ ),
    .B1(\MuI._1357_ ),
    .Y(\MuI._1358_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5560_  (.A(\MuI._1344_ ),
    .B(\MuI._1345_ ),
    .C(\MuI._1357_ ),
    .X(\MuI._1359_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5561_  (.A1(\MuI._1343_ ),
    .A2(\MuI._1358_ ),
    .B1_N(\MuI._1359_ ),
    .X(\MuI._1360_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5562_  (.A(\MuI._1313_ ),
    .B(\MuI._1317_ ),
    .C(\MuI._1319_ ),
    .X(\MuI._1361_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5563_  (.A1(\MuI._1313_ ),
    .A2(\MuI._1319_ ),
    .B1(\MuI._1317_ ),
    .Y(\MuI._1363_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5564_  (.A(\MuI._1361_ ),
    .B(\MuI._1363_ ),
    .Y(\MuI._1364_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5565_  (.A_N(\MuI._1360_ ),
    .B(\MuI._1364_ ),
    .X(\MuI._1365_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5566_  (.A(\MuI._1361_ ),
    .B(\MuI._1363_ ),
    .C(\MuI._1360_ ),
    .X(\MuI._1366_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5567_  (.A1(\MuI._1364_ ),
    .A2(\MuI._1359_ ),
    .B1(\MuI._1341_ ),
    .C1(\MuI._1366_ ),
    .X(\MuI._1367_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._5568_  (.A(\MuI._1323_ ),
    .B(\MuI._1324_ ),
    .C_N(\MuI._1325_ ),
    .X(\MuI._1368_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5569_  (.A1(\MuI._1323_ ),
    .A2(\MuI._1324_ ),
    .B1_N(\MuI._1325_ ),
    .Y(\MuI._1369_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5570_  (.A1(\MuI._1365_ ),
    .A2(\MuI._1367_ ),
    .B1(\MuI._1368_ ),
    .C1(\MuI._1369_ ),
    .Y(\MuI._1370_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5571_  (.A(\MuI._1334_ ),
    .B(\MuI._1370_ ),
    .Y(\MuI._1371_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5572_  (.A1(\MuI._1331_ ),
    .A2(\MuI._1332_ ),
    .B1(\MuI._1371_ ),
    .B2(\MuI._1294_ ),
    .X(\MuI._1372_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5573_  (.A1(\MuI._1368_ ),
    .A2(\MuI._1369_ ),
    .B1(\MuI._1365_ ),
    .C1(\MuI._1367_ ),
    .X(\MuI._1374_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5574_  (.A(\MuI._1364_ ),
    .B(\MuI._1360_ ),
    .Y(\MuI._1375_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._5575_  (.A(\MuI._1341_ ),
    .B(\MuI._1375_ ),
    .X(\MuI._1376_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5576_  (.A(\MuI._1356_ ),
    .B(\MuI._1347_ ),
    .C(\MuI._1355_ ),
    .Y(\MuI._1377_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5577_  (.A1(\MuI._1356_ ),
    .A2(\MuI._1355_ ),
    .B1(\MuI._1347_ ),
    .X(\MuI._1378_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5578_  (.A(\MuI._2886_ ),
    .B(\MuI._0245_ ),
    .Y(\MuI._1379_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5579_  (.A(\MuI._2882_ ),
    .B(\MuI._0320_ ),
    .Y(\MuI._1380_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5580_  (.A1(\MuI._2882_ ),
    .A2(\MuI._0315_ ),
    .B1(\MuI._0320_ ),
    .B2(\MuI._2886_ ),
    .X(\MuI._1381_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5581_  (.A1(\MuI._1379_ ),
    .A2(\MuI._1380_ ),
    .B1(\MuI._1381_ ),
    .X(\MuI._1382_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5582_  (.A(\MuI._1353_ ),
    .B(\MuI._1350_ ),
    .C(\MuI._1352_ ),
    .X(\MuI._1383_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5583_  (.A1(\MuI._1353_ ),
    .A2(\MuI._1352_ ),
    .B1(\MuI._1350_ ),
    .Y(\MuI._1385_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5584_  (.A(\MuI._3269_ ),
    .B(\MuI._0244_ ),
    .Y(\MuI._1386_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5585_  (.A1(\MuI._3397_ ),
    .A2(\MuI._0305_ ),
    .B1(\MuI._0111_ ),
    .B2(\MuI._3403_ ),
    .Y(\MuI._1387_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5586_  (.A(\MuI._3403_ ),
    .B(\MuI._3397_ ),
    .C(\MuI._3371_ ),
    .D(\MuI._0110_ ),
    .X(\MuI._1388_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5587_  (.A1(\MuI._1386_ ),
    .A2(\MuI._1387_ ),
    .B1_N(\MuI._1388_ ),
    .Y(\MuI._1389_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5588_  (.A1(\MuI._1383_ ),
    .A2(\MuI._1385_ ),
    .B1(\MuI._1389_ ),
    .X(\MuI._1390_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5589_  (.A(\MuI._1383_ ),
    .B(\MuI._1385_ ),
    .C(\MuI._1389_ ),
    .X(\MuI._1391_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5590_  (.A1(\MuI._1382_ ),
    .A2(\MuI._1390_ ),
    .B1(\MuI._1391_ ),
    .X(\MuI._1392_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5591_  (.A(\MuI._1377_ ),
    .B(\MuI._1378_ ),
    .C(\MuI._1392_ ),
    .X(\MuI._1393_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5592_  (.A1(\MuI._1377_ ),
    .A2(\MuI._1378_ ),
    .B1(\MuI._1392_ ),
    .Y(\MuI._1394_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5593_  (.A(\MuI._1379_ ),
    .B(\MuI._1380_ ),
    .Y(\MuI._1396_ ));
 sky130_fd_sc_hd__nor3b_1 \MuI._5594_  (.A(\MuI._1393_ ),
    .B(\MuI._1394_ ),
    .C_N(\MuI._1396_ ),
    .Y(\MuI._1397_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5595_  (.A(\MuI._1359_ ),
    .B(\MuI._1343_ ),
    .C(\MuI._1358_ ),
    .X(\MuI._1398_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5596_  (.A1(\MuI._1359_ ),
    .A2(\MuI._1358_ ),
    .B1(\MuI._1343_ ),
    .Y(\MuI._1399_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5597_  (.A1(\MuI._1393_ ),
    .A2(\MuI._1397_ ),
    .B1(\MuI._1398_ ),
    .C1(\MuI._1399_ ),
    .X(\MuI._1400_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5598_  (.A(\MuI._1370_ ),
    .B(\MuI._1374_ ),
    .C(\MuI._1376_ ),
    .D(\MuI._1400_ ),
    .Y(\MuI._1401_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5599_  (.A(\MuI._1334_ ),
    .B(\MuI._1401_ ),
    .X(\MuI._1402_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5600_  (.A1(\MuI._1365_ ),
    .A2(\MuI._1367_ ),
    .B1(\MuI._1368_ ),
    .C1(\MuI._1369_ ),
    .X(\MuI._1403_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5601_  (.A1(\MuI._1333_ ),
    .A2(\MuI._1403_ ),
    .B1(\MuI._1330_ ),
    .X(\MuI._1404_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5602_  (.A(\MuI._1292_ ),
    .B(\MuI._1293_ ),
    .C(\MuI._1404_ ),
    .X(\MuI._1405_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5603_  (.A1(\MuI._1292_ ),
    .A2(\MuI._1293_ ),
    .B1(\MuI._1404_ ),
    .Y(\MuI._1407_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5604_  (.A(\MuI._1402_ ),
    .B(\MuI._1405_ ),
    .C(\MuI._1407_ ),
    .Y(\MuI._1408_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5605_  (.A1(\MuI._1370_ ),
    .A2(\MuI._1374_ ),
    .B1(\MuI._1376_ ),
    .B2(\MuI._1400_ ),
    .X(\MuI._1409_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5606_  (.A1(\MuI._1398_ ),
    .A2(\MuI._1399_ ),
    .B1(\MuI._1393_ ),
    .C1(\MuI._1397_ ),
    .Y(\MuI._1410_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5607_  (.A1(\MuI._1393_ ),
    .A2(\MuI._1394_ ),
    .B1_N(\MuI._1396_ ),
    .X(\MuI._1411_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5608_  (.A(\MuI._1397_ ),
    .B(\MuI._1411_ ),
    .X(\MuI._1412_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5609_  (.A(\MuI._1412_ ),
    .Y(\MuI._1413_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5610_  (.A(\MuI._3397_ ),
    .B(\MuI._0245_ ),
    .X(\MuI._1414_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5611_  (.A(\MuI._3403_ ),
    .B(\MuI._0112_ ),
    .C(\MuI._1414_ ),
    .X(\MuI._1415_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5612_  (.A1(\MuI._3397_ ),
    .A2(\MuI._0112_ ),
    .B1(\MuI._0246_ ),
    .B2(\MuI._3403_ ),
    .Y(\MuI._1416_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._5613_  (.A_N(\MuI._1415_ ),
    .B_N(\MuI._1416_ ),
    .C(\MuI._3269_ ),
    .D(\MuI._0420_ ),
    .X(\MuI._1418_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5614_  (.A(\MuI._1388_ ),
    .B(\MuI._1387_ ),
    .Y(\MuI._1419_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5615_  (.A(\MuI._1386_ ),
    .B(\MuI._1419_ ),
    .Y(\MuI._1420_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5616_  (.A1(\MuI._1415_ ),
    .A2(\MuI._1418_ ),
    .B1(\MuI._1420_ ),
    .X(\MuI._1421_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5617_  (.A(\MuI._1420_ ),
    .B(\MuI._1415_ ),
    .C(\MuI._1418_ ),
    .Y(\MuI._1422_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5618_  (.A(\MuI._1380_ ),
    .B(\MuI._1421_ ),
    .C(\MuI._1422_ ),
    .Y(\MuI._1423_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5619_  (.A(\MuI._1391_ ),
    .B_N(\MuI._1390_ ),
    .X(\MuI._1424_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5620_  (.A(\MuI._1382_ ),
    .B(\MuI._1424_ ),
    .Y(\MuI._1425_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5621_  (.A1(\MuI._1421_ ),
    .A2(\MuI._1423_ ),
    .B1(\MuI._1425_ ),
    .X(\MuI._1426_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5622_  (.A(\MuI._1413_ ),
    .B(\MuI._1426_ ),
    .Y(\MuI._1427_ ));
 sky130_fd_sc_hd__or4b_1 \MuI._5623_  (.A(\MuI._1400_ ),
    .B(\MuI._1410_ ),
    .C(\MuI._1427_ ),
    .D_N(\MuI._1376_ ),
    .X(\MuI._1429_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5624_  (.A1(\MuI._1401_ ),
    .A2(\MuI._1409_ ),
    .B1_N(\MuI._1429_ ),
    .X(\MuI._1430_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5625_  (.A(\MuI._1400_ ),
    .B(\MuI._1410_ ),
    .Y(\MuI._1431_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5626_  (.A1(\MuI._1431_ ),
    .A2(\MuI._1413_ ),
    .A3(\MuI._1426_ ),
    .B1(\MuI._1400_ ),
    .X(\MuI._1432_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5627_  (.A(\MuI._1376_ ),
    .B(\MuI._1432_ ),
    .Y(\MuI._1433_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5628_  (.A(\MuI._1431_ ),
    .B(\MuI._1427_ ),
    .X(\MuI._1434_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5629_  (.A(\MuI._1425_ ),
    .B(\MuI._1421_ ),
    .C(\MuI._1423_ ),
    .Y(\MuI._1435_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5630_  (.A(\MuI._1426_ ),
    .B(\MuI._1435_ ),
    .Y(\MuI._1436_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5631_  (.A1(\MuI._1421_ ),
    .A2(\MuI._1422_ ),
    .B1(\MuI._1380_ ),
    .X(\MuI._1437_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5632_  (.A(\MuI._1423_ ),
    .B(\MuI._1437_ ),
    .Y(\MuI._1438_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5633_  (.A1_N(\MuI._3269_ ),
    .A2_N(\MuI._0421_ ),
    .B1(\MuI._1415_ ),
    .B2(\MuI._1416_ ),
    .X(\MuI._1440_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5634_  (.A(\MuI._1418_ ),
    .B(\MuI._1440_ ),
    .Y(\MuI._1441_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5635_  (.A(\MuI._3403_ ),
    .B(\MuI._0421_ ),
    .C(\MuI._1414_ ),
    .D(\MuI._1441_ ),
    .X(\MuI._1442_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5636_  (.A(\MuI._1438_ ),
    .B(\MuI._1442_ ),
    .X(\MuI._1443_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5637_  (.A(\MuI._1413_ ),
    .B(\MuI._1436_ ),
    .C(\MuI._1443_ ),
    .Y(\MuI._1444_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5638_  (.A(\MuI._1433_ ),
    .B(\MuI._1434_ ),
    .C(\MuI._1444_ ),
    .Y(\MuI._1445_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._5639_  (.A_N(\MuI._1429_ ),
    .B(\MuI._1409_ ),
    .C(\MuI._1401_ ),
    .X(\MuI._1446_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5640_  (.A1(\MuI._1430_ ),
    .A2(\MuI._1445_ ),
    .B1(\MuI._1446_ ),
    .X(\MuI._1447_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5641_  (.A(\MuI._1370_ ),
    .B(\MuI._1401_ ),
    .Y(\MuI._1448_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5642_  (.A(\MuI._1334_ ),
    .B(\MuI._1448_ ),
    .Y(\MuI._1449_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5643_  (.A1(\MuI._1405_ ),
    .A2(\MuI._1407_ ),
    .B1(\MuI._1402_ ),
    .Y(\MuI._1451_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5644_  (.A1(\MuI._1408_ ),
    .A2(\MuI._1447_ ),
    .A3(\MuI._1449_ ),
    .B1(\MuI._1451_ ),
    .X(\MuI._1452_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5645_  (.A(\MuI._1294_ ),
    .B(\MuI._1331_ ),
    .C(\MuI._1332_ ),
    .D(\MuI._1371_ ),
    .X(\MuI._1453_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5646_  (.A1(\MuI._1372_ ),
    .A2(\MuI._1452_ ),
    .B1(\MuI._1453_ ),
    .Y(\MuI._1454_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5647_  (.A(\MuI._1287_ ),
    .B(\MuI._1331_ ),
    .Y(\MuI._1455_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5648_  (.A(\MuI._1242_ ),
    .B(\MuI._1455_ ),
    .X(\MuI._1456_ ));
 sky130_fd_sc_hd__o22a_1 \MuI._5649_  (.A1(\MuI._1242_ ),
    .A2(\MuI._1331_ ),
    .B1(\MuI._1454_ ),
    .B2(\MuI._1456_ ),
    .X(\MuI._1457_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._5650_  (.A1(\MuI._1290_ ),
    .A2(\MuI._1457_ ),
    .B1(\MuI._1288_ ),
    .Y(\MuI._1458_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._5651_  (.A(\MuI._1062_ ),
    .B(\MuI._1172_ ),
    .C(\MuI._1178_ ),
    .Y(\MuI._1459_ ));
 sky130_fd_sc_hd__a221oi_4 \MuI._5652_  (.A1(\MuI._1182_ ),
    .A2(\MuI._1236_ ),
    .B1(\MuI._1239_ ),
    .B2(\MuI._1458_ ),
    .C1(\MuI._1459_ ),
    .Y(\MuI._1460_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5653_  (.A(\MuI._1062_ ),
    .B(\MuI._1179_ ),
    .Y(\MuI._1462_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5654_  (.A(\MuI._0984_ ),
    .B(\MuI._1060_ ),
    .Y(\MuI._1463_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._5655_  (.A1(\MuI._0844_ ),
    .A2(\MuI._1061_ ),
    .B1(\MuI._1463_ ),
    .X(\MuI._1464_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._5656_  (.A_N(\MuI._1057_ ),
    .B(\MuI._1058_ ),
    .C(\MuI._0992_ ),
    .X(\MuI._1465_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5657_  (.A(\MuI._1009_ ),
    .B(\MuI._1011_ ),
    .C(\MuI._1013_ ),
    .Y(\MuI._1466_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5658_  (.A1(\MuI._2860_ ),
    .A2(\MuI._0246_ ),
    .A3(\MuI._1005_ ),
    .B1(\MuI._1004_ ),
    .X(\MuI._1467_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5659_  (.A(\MuI._1318_ ),
    .B(\MuI._1813_ ),
    .C(\MuI._0246_ ),
    .D(\MuI._0420_ ),
    .Y(\MuI._1468_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5660_  (.A1(\MuI._1813_ ),
    .A2(\MuI._0246_ ),
    .B1(\MuI._0420_ ),
    .B2(\MuI._1318_ ),
    .X(\MuI._1469_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5661_  (.A(\MuI._1468_ ),
    .B(\MuI._1469_ ),
    .Y(\MuI._1470_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5662_  (.A(\MuI._1467_ ),
    .B(\MuI._1470_ ),
    .Y(\MuI._1471_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5663_  (.A(\MuI._0986_ ),
    .B(\MuI._1471_ ),
    .Y(\MuI._1473_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5664_  (.A(\MuI._0986_ ),
    .B(\MuI._1471_ ),
    .X(\MuI._1474_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5665_  (.A(\MuI._1473_ ),
    .B(\MuI._1474_ ),
    .Y(\MuI._1475_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5666_  (.A1(\MuI._1009_ ),
    .A2(\MuI._1466_ ),
    .B1(\MuI._1475_ ),
    .Y(\MuI._1476_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5667_  (.A(\MuI._1009_ ),
    .B(\MuI._1466_ ),
    .C(\MuI._1475_ ),
    .X(\MuI._1477_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5668_  (.A(\MuI._1476_ ),
    .B(\MuI._1477_ ),
    .Y(\MuI._1478_ ));
 sky130_fd_sc_hd__nor4_1 \MuI._5669_  (.A(\MuI._1014_ ),
    .B(\MuI._1015_ ),
    .C(\MuI._1052_ ),
    .D(\MuI._1053_ ),
    .Y(\MuI._1479_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5670_  (.A_N(\MuI._1001_ ),
    .B(\MuI._1000_ ),
    .X(\MuI._1480_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5671_  (.A(\MuI._1002_ ),
    .B(\MuI._1007_ ),
    .X(\MuI._1481_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5672_  (.A1(\MuI._1025_ ),
    .A2(\MuI._1026_ ),
    .B1_N(\MuI._1024_ ),
    .X(\MuI._1482_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5673_  (.A(\MuI.b_operand[11] ),
    .B(\MuI._2829_ ),
    .Y(\MuI._1484_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5674_  (.A(\MuI._2853_ ),
    .B(\MuI._2854_ ),
    .C(\MuI.a_operand[7] ),
    .D(\MuI.a_operand[6] ),
    .X(\MuI._1485_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5675_  (.A1(\MuI._2845_ ),
    .A2(\MuI._0088_ ),
    .B1(\MuI._2319_ ),
    .B2(\MuI._2844_ ),
    .Y(\MuI._1486_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5676_  (.A(\MuI._1484_ ),
    .B(\MuI._1485_ ),
    .C(\MuI._1486_ ),
    .X(\MuI._1487_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5677_  (.A1(\MuI._1485_ ),
    .A2(\MuI._1486_ ),
    .B1(\MuI._1484_ ),
    .Y(\MuI._1488_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5678_  (.A1(\MuI._2851_ ),
    .A2(\MuI._3247_ ),
    .A3(\MuI._0997_ ),
    .B1(\MuI._0996_ ),
    .X(\MuI._1489_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5679_  (.A(\MuI._1487_ ),
    .B(\MuI._1488_ ),
    .C(\MuI._1489_ ),
    .Y(\MuI._1490_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5680_  (.A1(\MuI._1487_ ),
    .A2(\MuI._1488_ ),
    .B1(\MuI._1489_ ),
    .X(\MuI._1491_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5681_  (.A(\MuI._2799_ ),
    .B(\MuI._2918_ ),
    .C(\MuI._0228_ ),
    .D(\MuI._3371_ ),
    .X(\MuI._1492_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5682_  (.A1(\MuI._2649_ ),
    .A2(\MuI._3246_ ),
    .B1(\MuI._0305_ ),
    .B2(\MuI._2704_ ),
    .Y(\MuI._1493_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5683_  (.A(\MuI._1492_ ),
    .B(\MuI._1493_ ),
    .X(\MuI._1495_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5684_  (.A(\MuI._2583_ ),
    .B(\MuI._0112_ ),
    .Y(\MuI._1496_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5685_  (.A(\MuI._1495_ ),
    .B(\MuI._1496_ ),
    .X(\MuI._1497_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5686_  (.A(\MuI._1490_ ),
    .B(\MuI._1491_ ),
    .C(\MuI._1497_ ),
    .Y(\MuI._1498_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5687_  (.A1(\MuI._1490_ ),
    .A2(\MuI._1491_ ),
    .B1(\MuI._1497_ ),
    .X(\MuI._1499_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5688_  (.A(\MuI._1482_ ),
    .B(\MuI._1498_ ),
    .C(\MuI._1499_ ),
    .Y(\MuI._1500_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5689_  (.A1(\MuI._1498_ ),
    .A2(\MuI._1499_ ),
    .B1(\MuI._1482_ ),
    .X(\MuI._1501_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5690_  (.A1(\MuI._1480_ ),
    .A2(\MuI._1481_ ),
    .B1(\MuI._1500_ ),
    .C1(\MuI._1501_ ),
    .Y(\MuI._1502_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5691_  (.A1(\MuI._1500_ ),
    .A2(\MuI._1501_ ),
    .B1(\MuI._1480_ ),
    .C1(\MuI._1481_ ),
    .X(\MuI._1503_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5692_  (.A(\MuI._1029_ ),
    .B(\MuI._1048_ ),
    .C(\MuI._1049_ ),
    .Y(\MuI._1504_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5693_  (.A1(\MuI._1033_ ),
    .A2(\MuI._1035_ ),
    .B1_N(\MuI._1031_ ),
    .Y(\MuI._1506_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5694_  (.A(\MuI._0168_ ),
    .B(\MuI._3349_ ),
    .Y(\MuI._1507_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5695_  (.A(\MuI._2790_ ),
    .B(\MuI._2867_ ),
    .C(\MuI._3223_ ),
    .D(\MuI._2875_ ),
    .Y(\MuI._1508_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5696_  (.A1(\MuI._2873_ ),
    .A2(\MuI._2785_ ),
    .B1(\MuI._2875_ ),
    .B2(\MuI._2765_ ),
    .X(\MuI._1509_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._5697_  (.A_N(\MuI._1507_ ),
    .B(\MuI._1508_ ),
    .C(\MuI._1509_ ),
    .Y(\MuI._1510_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5698_  (.A1(\MuI._1508_ ),
    .A2(\MuI._1509_ ),
    .B1_N(\MuI._1507_ ),
    .X(\MuI._1511_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5699_  (.A(\MuI._1506_ ),
    .B(\MuI._1510_ ),
    .C(\MuI._1511_ ),
    .X(\MuI._1512_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5700_  (.A1(\MuI._1510_ ),
    .A2(\MuI._1511_ ),
    .B1(\MuI._1506_ ),
    .Y(\MuI._1513_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5701_  (.A(\MuI._1019_ ),
    .B(\MuI._1022_ ),
    .X(\MuI._1514_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5702_  (.A(\MuI._1512_ ),
    .B(\MuI._1513_ ),
    .C(\MuI._1514_ ),
    .X(\MuI._1515_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5703_  (.A1(\MuI._1512_ ),
    .A2(\MuI._1513_ ),
    .B1(\MuI._1514_ ),
    .Y(\MuI._1517_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5704_  (.A(\MuI._1515_ ),
    .B(\MuI._1517_ ),
    .X(\MuI._1518_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5705_  (.A1(\MuI._1036_ ),
    .A2(\MuI._1045_ ),
    .B1_N(\MuI._1044_ ),
    .X(\MuI._1519_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5706_  (.A1(\MuI._2451_ ),
    .A2(\MuI._2892_ ),
    .B1(\MuI._3185_ ),
    .B2(\MuI._2440_ ),
    .Y(\MuI._1520_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5707_  (.A(\MuI._2429_ ),
    .B(\MuI._0327_ ),
    .C(\MuI._2885_ ),
    .D(\MuI._3307_ ),
    .X(\MuI._1521_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5708_  (.A(\MuI._1520_ ),
    .B(\MuI._1521_ ),
    .Y(\MuI._1522_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5709_  (.A(\MuI._2484_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._1523_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5710_  (.A(\MuI._1522_ ),
    .B(\MuI._1523_ ),
    .Y(\MuI._1524_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5711_  (.A1(\MuI._1038_ ),
    .A2(\MuI._1040_ ),
    .B1_N(\MuI._1039_ ),
    .Y(\MuI._1525_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5712_  (.A(\MuI._2660_ ),
    .B(\MuI._0378_ ),
    .Y(\MuI._1526_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5713_  (.A(\MuI._2852_ ),
    .B(\MuI.a_operand[15] ),
    .C(\MuI._0017_ ),
    .D(\MuI._3396_ ),
    .X(\MuI._1528_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._5714_  (.A1(\MuI._2605_ ),
    .A2(\MuI._3262_ ),
    .B1(\MuI._0020_ ),
    .B2(\MuI._2852_ ),
    .Y(\MuI._1529_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5715_  (.A(\MuI._1526_ ),
    .B(\MuI._1528_ ),
    .C(\MuI._1529_ ),
    .X(\MuI._1530_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5716_  (.A1(\MuI._1528_ ),
    .A2(\MuI._1529_ ),
    .B1(\MuI._1526_ ),
    .Y(\MuI._1531_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5717_  (.A(\MuI._1525_ ),
    .B(\MuI._1530_ ),
    .C(\MuI._1531_ ),
    .Y(\MuI._1532_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5718_  (.A1(\MuI._1530_ ),
    .A2(\MuI._1531_ ),
    .B1(\MuI._1525_ ),
    .X(\MuI._1533_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5719_  (.A(\MuI._1524_ ),
    .B(\MuI._1532_ ),
    .C(\MuI._1533_ ),
    .Y(\MuI._1534_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5720_  (.A1(\MuI._1532_ ),
    .A2(\MuI._1533_ ),
    .B1(\MuI._1524_ ),
    .X(\MuI._1535_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._5721_  (.A(\MuI._1519_ ),
    .B(\MuI._1534_ ),
    .C(\MuI._1535_ ),
    .Y(\MuI._1536_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5722_  (.A1(\MuI._1534_ ),
    .A2(\MuI._1535_ ),
    .B1(\MuI._1519_ ),
    .X(\MuI._1537_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5723_  (.A(\MuI._1518_ ),
    .B(\MuI._1536_ ),
    .C(\MuI._1537_ ),
    .X(\MuI._1539_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5724_  (.A1(\MuI._1536_ ),
    .A2(\MuI._1537_ ),
    .B1(\MuI._1518_ ),
    .Y(\MuI._1540_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5725_  (.A1(\MuI._1048_ ),
    .A2(\MuI._1504_ ),
    .B1(\MuI._1539_ ),
    .C1(\MuI._1540_ ),
    .X(\MuI._1541_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5726_  (.A1(\MuI._1539_ ),
    .A2(\MuI._1540_ ),
    .B1(\MuI._1048_ ),
    .C1(\MuI._1504_ ),
    .Y(\MuI._1542_ ));
 sky130_fd_sc_hd__nand4_2 \MuI._5727_  (.A(\MuI._1502_ ),
    .B(\MuI._1503_ ),
    .C(\MuI._1541_ ),
    .D(\MuI._1542_ ),
    .Y(\MuI._1543_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5728_  (.A1(\MuI._1502_ ),
    .A2(\MuI._1503_ ),
    .B1(\MuI._1541_ ),
    .B2(\MuI._1542_ ),
    .X(\MuI._1544_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._5729_  (.A1(\MuI._1052_ ),
    .A2(\MuI._1479_ ),
    .B1(\MuI._1543_ ),
    .C1(\MuI._1544_ ),
    .Y(\MuI._1545_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5730_  (.A1(\MuI._1543_ ),
    .A2(\MuI._1544_ ),
    .B1(\MuI._1052_ ),
    .C1(\MuI._1479_ ),
    .X(\MuI._1546_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5731_  (.A(\MuI._1478_ ),
    .B(\MuI._1545_ ),
    .C(\MuI._1546_ ),
    .Y(\MuI._1547_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5732_  (.A1(\MuI._1545_ ),
    .A2(\MuI._1546_ ),
    .B1(\MuI._1478_ ),
    .X(\MuI._1548_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5733_  (.A1(\MuI._1057_ ),
    .A2(\MuI._1465_ ),
    .B1(\MuI._1547_ ),
    .C1(\MuI._1548_ ),
    .Y(\MuI._1550_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5734_  (.A1(\MuI._1547_ ),
    .A2(\MuI._1548_ ),
    .B1(\MuI._1057_ ),
    .C1(\MuI._1465_ ),
    .X(\MuI._1551_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5735_  (.A(\MuI._0990_ ),
    .B(\MuI._1550_ ),
    .C(\MuI._1551_ ),
    .X(\MuI._1552_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5736_  (.A1(\MuI._1550_ ),
    .A2(\MuI._1551_ ),
    .B1(\MuI._0990_ ),
    .Y(\MuI._1553_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5737_  (.A(\MuI._1552_ ),
    .B(\MuI._1553_ ),
    .Y(\MuI._1554_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5738_  (.A(\MuI._1464_ ),
    .B(\MuI._1554_ ),
    .Y(\MuI._1555_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5739_  (.A(\MuI._1464_ ),
    .B(\MuI._1552_ ),
    .C(\MuI._1553_ ),
    .X(\MuI._1556_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5740_  (.A1(\MuI._0990_ ),
    .A2(\MuI._1551_ ),
    .B1_N(\MuI._1550_ ),
    .X(\MuI._1557_ ));
 sky130_fd_sc_hd__o21bai_2 \MuI._5741_  (.A1(\MuI._1495_ ),
    .A2(\MuI._1496_ ),
    .B1_N(\MuI._1492_ ),
    .Y(\MuI._1558_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5742_  (.A(\MuI._1274_ ),
    .B(\MuI._0320_ ),
    .Y(\MuI._1559_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5743_  (.A(\MuI._3000_ ),
    .B(\MuI._2754_ ),
    .C(\MuI._0110_ ),
    .D(\MuI.a_operand[1] ),
    .X(\MuI._1561_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5744_  (.A1(\MuI._2754_ ),
    .A2(\MuI._0110_ ),
    .B1(\MuI.a_operand[1] ),
    .B2(\MuI._1307_ ),
    .X(\MuI._1562_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5745_  (.A_N(\MuI._1561_ ),
    .B(\MuI._1562_ ),
    .X(\MuI._1563_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5746_  (.A(\MuI._1559_ ),
    .B(\MuI._1563_ ),
    .Y(\MuI._1564_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5747_  (.A(\MuI._1558_ ),
    .B(\MuI._1564_ ),
    .Y(\MuI._1565_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5748_  (.A(\MuI._1318_ ),
    .B(\MuI._1813_ ),
    .C(\MuI._0245_ ),
    .D(\MuI._0320_ ),
    .X(\MuI._1566_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5749_  (.A1(\MuI._1467_ ),
    .A2(\MuI._1469_ ),
    .B1(\MuI._1566_ ),
    .Y(\MuI._1567_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5750_  (.A(\MuI._1565_ ),
    .B(\MuI._1567_ ),
    .Y(\MuI._1568_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5751_  (.A1(\MuI._1500_ ),
    .A2(\MuI._1502_ ),
    .B1(\MuI._1568_ ),
    .X(\MuI._1569_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5752_  (.A(\MuI._1500_ ),
    .B(\MuI._1502_ ),
    .C(\MuI._1568_ ),
    .Y(\MuI._1570_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5753_  (.A(\MuI._1569_ ),
    .B(\MuI._1570_ ),
    .Y(\MuI._1572_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5754_  (.A(\MuI._1473_ ),
    .B(\MuI._1572_ ),
    .X(\MuI._1573_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5755_  (.A1(\MuI._1513_ ),
    .A2(\MuI._1514_ ),
    .B1_N(\MuI._1512_ ),
    .Y(\MuI._1574_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5756_  (.A(\MuI.b_operand[11] ),
    .B(\MuI._3362_ ),
    .Y(\MuI._1575_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._5757_  (.A(\MuI._2836_ ),
    .B(\MuI._2838_ ),
    .C(\MuI._3349_ ),
    .D(\MuI._0085_ ),
    .Y(\MuI._1576_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5758_  (.A1(\MuI._2854_ ),
    .A2(\MuI._2341_ ),
    .B1(\MuI._0085_ ),
    .B2(\MuI._2853_ ),
    .X(\MuI._1577_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._5759_  (.A_N(\MuI._1575_ ),
    .B(\MuI._1576_ ),
    .C(\MuI._1577_ ),
    .Y(\MuI._1578_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5760_  (.A1(\MuI._1576_ ),
    .A2(\MuI._1577_ ),
    .B1_N(\MuI._1575_ ),
    .X(\MuI._1579_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5761_  (.A1(\MuI._1484_ ),
    .A2(\MuI._1486_ ),
    .B1_N(\MuI._1485_ ),
    .Y(\MuI._1580_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5762_  (.A(\MuI._1578_ ),
    .B(\MuI._1579_ ),
    .C(\MuI._1580_ ),
    .X(\MuI._1581_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5763_  (.A1(\MuI._1578_ ),
    .A2(\MuI._1579_ ),
    .B1(\MuI._1580_ ),
    .Y(\MuI._1583_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5764_  (.A(\MuI._2796_ ),
    .B(\MuI._0305_ ),
    .Y(\MuI._1584_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5765_  (.A(\MuI._2693_ ),
    .B(\MuI._2638_ ),
    .C(\MuI._2829_ ),
    .D(\MuI._3245_ ),
    .X(\MuI._1585_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5766_  (.A1(\MuI._2803_ ),
    .A2(\MuI._2829_ ),
    .B1(\MuI._3246_ ),
    .B2(\MuI._2802_ ),
    .Y(\MuI._1586_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5767_  (.A(\MuI._1585_ ),
    .B(\MuI._1586_ ),
    .Y(\MuI._1587_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5768_  (.A(\MuI._1584_ ),
    .B(\MuI._1587_ ),
    .Y(\MuI._1588_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._5769_  (.A(\MuI._1581_ ),
    .B(\MuI._1583_ ),
    .C_N(\MuI._1588_ ),
    .X(\MuI._1589_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5770_  (.A1(\MuI._1581_ ),
    .A2(\MuI._1583_ ),
    .B1_N(\MuI._1588_ ),
    .Y(\MuI._1590_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5771_  (.A(\MuI._1574_ ),
    .B(\MuI._1589_ ),
    .C(\MuI._1590_ ),
    .Y(\MuI._1591_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5772_  (.A1(\MuI._1589_ ),
    .A2(\MuI._1590_ ),
    .B1(\MuI._1574_ ),
    .X(\MuI._1592_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5773_  (.A(\MuI._1490_ ),
    .B(\MuI._1498_ ),
    .Y(\MuI._1594_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5774_  (.A(\MuI._1591_ ),
    .B(\MuI._1592_ ),
    .C(\MuI._1594_ ),
    .X(\MuI._1595_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5775_  (.A1(\MuI._1591_ ),
    .A2(\MuI._1592_ ),
    .B1(\MuI._1594_ ),
    .Y(\MuI._1596_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5776_  (.A(\MuI._1518_ ),
    .B(\MuI._1536_ ),
    .C(\MuI._1537_ ),
    .Y(\MuI._1597_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5777_  (.A1(\MuI._1520_ ),
    .A2(\MuI._1523_ ),
    .B1_N(\MuI._1521_ ),
    .X(\MuI._1598_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5778_  (.A(\MuI._0168_ ),
    .B(\MuI._3223_ ),
    .Y(\MuI._1599_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5779_  (.A(\MuI._0477_ ),
    .B(\MuI.a_operand[10] ),
    .C(\MuI._2866_ ),
    .D(\MuI._2868_ ),
    .X(\MuI._1600_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5780_  (.A1(\MuI._2765_ ),
    .A2(\MuI._3189_ ),
    .B1(\MuI._2875_ ),
    .B2(\MuI._0477_ ),
    .Y(\MuI._1601_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5781_  (.A(\MuI._1600_ ),
    .B(\MuI._1601_ ),
    .Y(\MuI._1602_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5782_  (.A(\MuI._1599_ ),
    .B(\MuI._1602_ ),
    .Y(\MuI._1603_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5783_  (.A(\MuI._1598_ ),
    .B(\MuI._1603_ ),
    .Y(\MuI._1605_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5784_  (.A(\MuI._1508_ ),
    .B(\MuI._1510_ ),
    .X(\MuI._1606_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5785_  (.A(\MuI._1605_ ),
    .B(\MuI._1606_ ),
    .Y(\MuI._1607_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5786_  (.A1(\MuI._1524_ ),
    .A2(\MuI._1533_ ),
    .B1_N(\MuI._1532_ ),
    .X(\MuI._1608_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5787_  (.A(\MuI._0743_ ),
    .B(\MuI._0741_ ),
    .C(\MuI._0742_ ),
    .X(\MuI._1609_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._5788_  (.A1(\MuI._1526_ ),
    .A2(\MuI._1529_ ),
    .B1_N(\MuI._1528_ ),
    .Y(\MuI._1610_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5789_  (.A1(\MuI._0743_ ),
    .A2(\MuI._0742_ ),
    .B1(\MuI._0741_ ),
    .Y(\MuI._1611_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5790_  (.A(\MuI._1609_ ),
    .B(\MuI._1610_ ),
    .C(\MuI._1611_ ),
    .Y(\MuI._1612_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5791_  (.A1(\MuI._1609_ ),
    .A2(\MuI._1611_ ),
    .B1(\MuI._1610_ ),
    .X(\MuI._1613_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5792_  (.A(\MuI._2451_ ),
    .B(\MuI._2966_ ),
    .Y(\MuI._1614_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._5793_  (.A1(\MuI._2429_ ),
    .A2(\MuI._3306_ ),
    .B1(\MuI._2881_ ),
    .B2(\MuI._2660_ ),
    .Y(\MuI._1616_ ));
 sky130_fd_sc_hd__and4_1 \MuI._5794_  (.A(\MuI._2660_ ),
    .B(\MuI._2429_ ),
    .C(\MuI._3306_ ),
    .D(\MuI._2880_ ),
    .X(\MuI._1617_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5795_  (.A(\MuI._1616_ ),
    .B(\MuI._1617_ ),
    .Y(\MuI._1618_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5796_  (.A(\MuI._1614_ ),
    .B(\MuI._1618_ ),
    .Y(\MuI._1619_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5797_  (.A(\MuI._1612_ ),
    .B(\MuI._1613_ ),
    .C(\MuI._1619_ ),
    .Y(\MuI._1620_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5798_  (.A1(\MuI._1612_ ),
    .A2(\MuI._1613_ ),
    .B1(\MuI._1619_ ),
    .X(\MuI._1621_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5799_  (.A(\MuI._1608_ ),
    .B(\MuI._1620_ ),
    .C(\MuI._1621_ ),
    .Y(\MuI._1622_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5800_  (.A1(\MuI._1620_ ),
    .A2(\MuI._1621_ ),
    .B1(\MuI._1608_ ),
    .X(\MuI._1623_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5801_  (.A(\MuI._1607_ ),
    .B(\MuI._1622_ ),
    .C(\MuI._1623_ ),
    .X(\MuI._1624_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5802_  (.A1(\MuI._1622_ ),
    .A2(\MuI._1623_ ),
    .B1(\MuI._1607_ ),
    .Y(\MuI._1625_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._5803_  (.A1(\MuI._1536_ ),
    .A2(\MuI._1597_ ),
    .B1(\MuI._1624_ ),
    .C1(\MuI._1625_ ),
    .Y(\MuI._1627_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5804_  (.A1(\MuI._1624_ ),
    .A2(\MuI._1625_ ),
    .B1(\MuI._1536_ ),
    .C1(\MuI._1597_ ),
    .X(\MuI._1628_ ));
 sky130_fd_sc_hd__nor4_2 \MuI._5805_  (.A(\MuI._1595_ ),
    .B(\MuI._1596_ ),
    .C(\MuI._1627_ ),
    .D(\MuI._1628_ ),
    .Y(\MuI._1629_ ));
 sky130_fd_sc_hd__o22a_1 \MuI._5806_  (.A1(\MuI._1595_ ),
    .A2(\MuI._1596_ ),
    .B1(\MuI._1627_ ),
    .B2(\MuI._1628_ ),
    .X(\MuI._1630_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5807_  (.A1(\MuI._1541_ ),
    .A2(\MuI._1543_ ),
    .B1(\MuI._1629_ ),
    .C1(\MuI._1630_ ),
    .X(\MuI._1631_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5808_  (.A1(\MuI._1629_ ),
    .A2(\MuI._1630_ ),
    .B1(\MuI._1541_ ),
    .C1(\MuI._1543_ ),
    .Y(\MuI._1632_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5809_  (.A(\MuI._1573_ ),
    .B(\MuI._1631_ ),
    .C(\MuI._1632_ ),
    .X(\MuI._1633_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5810_  (.A1(\MuI._1631_ ),
    .A2(\MuI._1632_ ),
    .B1(\MuI._1573_ ),
    .Y(\MuI._1634_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5811_  (.A1(\MuI._1545_ ),
    .A2(\MuI._1547_ ),
    .B1(\MuI._1633_ ),
    .C1(\MuI._1634_ ),
    .X(\MuI._1635_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5812_  (.A1(\MuI._1633_ ),
    .A2(\MuI._1634_ ),
    .B1(\MuI._1545_ ),
    .C1(\MuI._1547_ ),
    .Y(\MuI._1636_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5813_  (.A(\MuI._1476_ ),
    .B(\MuI._1635_ ),
    .C(\MuI._1636_ ),
    .X(\MuI._1638_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5814_  (.A1(\MuI._1635_ ),
    .A2(\MuI._1636_ ),
    .B1(\MuI._1476_ ),
    .Y(\MuI._1639_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5815_  (.A(\MuI._1638_ ),
    .B(\MuI._1639_ ),
    .Y(\MuI._1640_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5816_  (.A(\MuI._1557_ ),
    .B(\MuI._1640_ ),
    .Y(\MuI._1641_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5817_  (.A(\MuI._1556_ ),
    .B(\MuI._1641_ ),
    .Y(\MuI._1642_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5818_  (.A(\MuI._1462_ ),
    .B(\MuI._1555_ ),
    .Y(\MuI._1643_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5819_  (.A_N(\MuI._1642_ ),
    .B(\MuI._1643_ ),
    .X(\MuI._1644_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5820_  (.A1(\MuI._1462_ ),
    .A2(\MuI._1555_ ),
    .B1(\MuI._1644_ ),
    .Y(\MuI._1645_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5821_  (.A(\MuI._1557_ ),
    .B(\MuI._1640_ ),
    .Y(\MuI._1646_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5822_  (.A1(\MuI._1476_ ),
    .A2(\MuI._1636_ ),
    .B1_N(\MuI._1635_ ),
    .X(\MuI._1647_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5823_  (.A1(\MuI._1473_ ),
    .A2(\MuI._1572_ ),
    .B1(\MuI._1569_ ),
    .Y(\MuI._1649_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5824_  (.A(\MuI._1573_ ),
    .B(\MuI._1631_ ),
    .C(\MuI._1632_ ),
    .Y(\MuI._1650_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5825_  (.A1(\MuI._1574_ ),
    .A2(\MuI._1589_ ),
    .A3(\MuI._1590_ ),
    .B1(\MuI._1595_ ),
    .X(\MuI._1651_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5826_  (.A(\MuI._1164_ ),
    .B(\MuI._0421_ ),
    .Y(\MuI._1652_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5827_  (.A1(\MuI._1285_ ),
    .A2(\MuI._0321_ ),
    .A3(\MuI._1562_ ),
    .B1(\MuI._1561_ ),
    .X(\MuI._1653_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5828_  (.A1(\MuI._1584_ ),
    .A2(\MuI._1586_ ),
    .B1_N(\MuI._1585_ ),
    .X(\MuI._1654_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5829_  (.A(\MuI._1263_ ),
    .B(\MuI._0244_ ),
    .Y(\MuI._1655_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5830_  (.A_N(\MuI._0718_ ),
    .B(\MuI._0717_ ),
    .X(\MuI._1656_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5831_  (.A(\MuI._1655_ ),
    .B(\MuI._1656_ ),
    .Y(\MuI._1657_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5832_  (.A(\MuI._1654_ ),
    .B(\MuI._1657_ ),
    .Y(\MuI._1658_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._5833_  (.A(\MuI._1653_ ),
    .B(\MuI._1658_ ),
    .Y(\MuI._1660_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5834_  (.A1(\MuI._1558_ ),
    .A2(\MuI._1564_ ),
    .B1(\MuI._1566_ ),
    .X(\MuI._1661_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._5835_  (.A1(\MuI._1558_ ),
    .A2(\MuI._1564_ ),
    .B1(\MuI._1661_ ),
    .Y(\MuI._1662_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5836_  (.A(\MuI._1660_ ),
    .B(\MuI._1662_ ),
    .X(\MuI._1663_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5837_  (.A(\MuI._1652_ ),
    .B(\MuI._1663_ ),
    .Y(\MuI._1664_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5838_  (.A(\MuI._1651_ ),
    .B(\MuI._1664_ ),
    .Y(\MuI._1665_ ));
 sky130_fd_sc_hd__and4b_1 \MuI._5839_  (.A_N(\MuI._1565_ ),
    .B(\MuI._1469_ ),
    .C(\MuI._1468_ ),
    .D(\MuI._1467_ ),
    .X(\MuI._1666_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5840_  (.A(\MuI._1665_ ),
    .B(\MuI._1666_ ),
    .Y(\MuI._1667_ ));
 sky130_fd_sc_hd__nor3b_1 \MuI._5841_  (.A(\MuI._1581_ ),
    .B(\MuI._1583_ ),
    .C_N(\MuI._1588_ ),
    .Y(\MuI._1668_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5842_  (.A(\MuI._1598_ ),
    .B_N(\MuI._1603_ ),
    .X(\MuI._1669_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5843_  (.A(\MuI._1606_ ),
    .B_N(\MuI._1605_ ),
    .X(\MuI._1671_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5844_  (.A1_N(\MuI.b_operand[11] ),
    .A2_N(\MuI._0088_ ),
    .B1(\MuI._0694_ ),
    .B2(\MuI._0695_ ),
    .X(\MuI._1672_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5845_  (.A(\MuI._0696_ ),
    .B(\MuI._1672_ ),
    .Y(\MuI._1673_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5846_  (.A(\MuI._1576_ ),
    .B(\MuI._1578_ ),
    .Y(\MuI._1674_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5847_  (.A(\MuI._1673_ ),
    .B(\MuI._1674_ ),
    .X(\MuI._1675_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5848_  (.A1_N(\MuI._2796_ ),
    .A2_N(\MuI._3247_ ),
    .B1(\MuI._0710_ ),
    .B2(\MuI._0711_ ),
    .X(\MuI._1676_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5849_  (.A(\MuI._0712_ ),
    .B(\MuI._1676_ ),
    .Y(\MuI._1677_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5850_  (.A(\MuI._1675_ ),
    .B(\MuI._1677_ ),
    .Y(\MuI._1678_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5851_  (.A1(\MuI._1669_ ),
    .A2(\MuI._1671_ ),
    .B1(\MuI._1678_ ),
    .X(\MuI._1679_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5852_  (.A(\MuI._1669_ ),
    .B(\MuI._1671_ ),
    .C(\MuI._1678_ ),
    .Y(\MuI._1680_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5853_  (.A1(\MuI._1581_ ),
    .A2(\MuI._1668_ ),
    .B1(\MuI._1679_ ),
    .C1(\MuI._1680_ ),
    .X(\MuI._1682_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5854_  (.A1(\MuI._1679_ ),
    .A2(\MuI._1680_ ),
    .B1(\MuI._1581_ ),
    .C1(\MuI._1668_ ),
    .Y(\MuI._1683_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5855_  (.A(\MuI._1607_ ),
    .B(\MuI._1622_ ),
    .C(\MuI._1623_ ),
    .Y(\MuI._1684_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5856_  (.A1(\MuI._1613_ ),
    .A2(\MuI._1619_ ),
    .B1_N(\MuI._1612_ ),
    .X(\MuI._1685_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5857_  (.A1(\MuI._0747_ ),
    .A2(\MuI._0748_ ),
    .B1(\MuI._0749_ ),
    .X(\MuI._1686_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5858_  (.A(\MuI._0750_ ),
    .B(\MuI._1685_ ),
    .C(\MuI._1686_ ),
    .Y(\MuI._1687_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5859_  (.A1(\MuI._0750_ ),
    .A2(\MuI._1686_ ),
    .B1(\MuI._1685_ ),
    .X(\MuI._1688_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5860_  (.A1(\MuI._1599_ ),
    .A2(\MuI._1601_ ),
    .B1_N(\MuI._1600_ ),
    .X(\MuI._1689_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._5861_  (.A1(\MuI._1614_ ),
    .A2(\MuI._1616_ ),
    .B1_N(\MuI._1617_ ),
    .X(\MuI._1690_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._5862_  (.A1_N(\MuI._2790_ ),
    .A2_N(\MuI._0168_ ),
    .B1(\MuI._0683_ ),
    .B2(\MuI._0684_ ),
    .X(\MuI._1691_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5863_  (.A(\MuI._0685_ ),
    .B(\MuI._1691_ ),
    .Y(\MuI._1693_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5864_  (.A(\MuI._1690_ ),
    .B(\MuI._1693_ ),
    .Y(\MuI._1694_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5865_  (.A(\MuI._1689_ ),
    .B(\MuI._1694_ ),
    .Y(\MuI._1695_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5866_  (.A(\MuI._1687_ ),
    .B(\MuI._1688_ ),
    .C(\MuI._1695_ ),
    .X(\MuI._1696_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5867_  (.A1(\MuI._1687_ ),
    .A2(\MuI._1688_ ),
    .B1(\MuI._1695_ ),
    .Y(\MuI._1697_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5868_  (.A1(\MuI._1622_ ),
    .A2(\MuI._1684_ ),
    .B1(\MuI._1696_ ),
    .C1(\MuI._1697_ ),
    .Y(\MuI._1698_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5869_  (.A1(\MuI._1696_ ),
    .A2(\MuI._1697_ ),
    .B1(\MuI._1622_ ),
    .C1(\MuI._1684_ ),
    .X(\MuI._1699_ ));
 sky130_fd_sc_hd__or4_1 \MuI._5870_  (.A(\MuI._1682_ ),
    .B(\MuI._1683_ ),
    .C(\MuI._1698_ ),
    .D(\MuI._1699_ ),
    .X(\MuI._1700_ ));
 sky130_fd_sc_hd__o22ai_1 \MuI._5871_  (.A1(\MuI._1682_ ),
    .A2(\MuI._1683_ ),
    .B1(\MuI._1698_ ),
    .B2(\MuI._1699_ ),
    .Y(\MuI._1701_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5872_  (.A1(\MuI._1627_ ),
    .A2(\MuI._1629_ ),
    .B1(\MuI._1700_ ),
    .C1(\MuI._1701_ ),
    .Y(\MuI._1702_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5873_  (.A1(\MuI._1700_ ),
    .A2(\MuI._1701_ ),
    .B1(\MuI._1627_ ),
    .C1(\MuI._1629_ ),
    .X(\MuI._1704_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5874_  (.A(\MuI._1667_ ),
    .B(\MuI._1702_ ),
    .C(\MuI._1704_ ),
    .X(\MuI._1705_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5875_  (.A1(\MuI._1702_ ),
    .A2(\MuI._1704_ ),
    .B1(\MuI._1667_ ),
    .Y(\MuI._1706_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5876_  (.A1(\MuI._1631_ ),
    .A2(\MuI._1650_ ),
    .B1(\MuI._1705_ ),
    .C1(\MuI._1706_ ),
    .X(\MuI._1707_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5877_  (.A1(\MuI._1705_ ),
    .A2(\MuI._1706_ ),
    .B1(\MuI._1631_ ),
    .C1(\MuI._1650_ ),
    .Y(\MuI._1708_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5878_  (.A(\MuI._1707_ ),
    .B(\MuI._1708_ ),
    .Y(\MuI._1709_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5879_  (.A(\MuI._1649_ ),
    .B(\MuI._1709_ ),
    .Y(\MuI._1710_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5880_  (.A(\MuI._1647_ ),
    .B(\MuI._1710_ ),
    .Y(\MuI._1711_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5881_  (.A(\MuI._1646_ ),
    .B(\MuI._1711_ ),
    .Y(\MuI._1712_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5882_  (.A(\MuI._1647_ ),
    .B(\MuI._1710_ ),
    .Y(\MuI._1713_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5883_  (.A_N(\MuI._1665_ ),
    .B(\MuI._1666_ ),
    .X(\MuI._1715_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5884_  (.A1(\MuI._1651_ ),
    .A2(\MuI._1664_ ),
    .B1(\MuI._1715_ ),
    .X(\MuI._1716_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._5885_  (.A1(\MuI._1667_ ),
    .A2(\MuI._1704_ ),
    .B1_N(\MuI._1702_ ),
    .Y(\MuI._1717_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5886_  (.A(\MuI._1660_ ),
    .B(\MuI._1662_ ),
    .Y(\MuI._1718_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5887_  (.A(\MuI._1164_ ),
    .B(\MuI._0421_ ),
    .C(\MuI._1663_ ),
    .X(\MuI._1719_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5888_  (.A1(\MuI._1581_ ),
    .A2(\MuI._1668_ ),
    .B1(\MuI._1679_ ),
    .C1(\MuI._1680_ ),
    .Y(\MuI._1720_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5889_  (.A(\MuI._1654_ ),
    .B_N(\MuI._1657_ ),
    .X(\MuI._1721_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5890_  (.A(\MuI._1653_ ),
    .B(\MuI._1658_ ),
    .Y(\MuI._1722_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5891_  (.A(\MuI._0719_ ),
    .B(\MuI._0721_ ),
    .Y(\MuI._1723_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._5892_  (.A1(\MuI._1721_ ),
    .A2(\MuI._1722_ ),
    .B1(\MuI._1723_ ),
    .Y(\MuI._1724_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5893_  (.A(\MuI._1721_ ),
    .B(\MuI._1722_ ),
    .C(\MuI._1723_ ),
    .X(\MuI._1726_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._5894_  (.A1(\MuI._1164_ ),
    .A2(\MuI._0246_ ),
    .B1(\MuI._0420_ ),
    .B2(\MuI._0746_ ),
    .X(\MuI._1727_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5895_  (.A(\MuI._1727_ ),
    .Y(\MuI._1728_ ));
 sky130_fd_sc_hd__nor4_1 \MuI._5896_  (.A(\MuI._0727_ ),
    .B(\MuI._1724_ ),
    .C(\MuI._1726_ ),
    .D(\MuI._1728_ ),
    .Y(\MuI._1729_ ));
 sky130_fd_sc_hd__o22a_1 \MuI._5897_  (.A1(\MuI._1724_ ),
    .A2(\MuI._1726_ ),
    .B1(\MuI._1728_ ),
    .B2(\MuI._0727_ ),
    .X(\MuI._1730_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5898_  (.A1(\MuI._1679_ ),
    .A2(\MuI._1720_ ),
    .B1(\MuI._1729_ ),
    .C1(\MuI._1730_ ),
    .X(\MuI._1731_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5899_  (.A1(\MuI._1729_ ),
    .A2(\MuI._1730_ ),
    .B1(\MuI._1679_ ),
    .C1(\MuI._1720_ ),
    .Y(\MuI._1732_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5900_  (.A1(\MuI._1718_ ),
    .A2(\MuI._1719_ ),
    .B1(\MuI._1731_ ),
    .C1(\MuI._1732_ ),
    .Y(\MuI._1733_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5901_  (.A1(\MuI._1731_ ),
    .A2(\MuI._1732_ ),
    .B1(\MuI._1718_ ),
    .C1(\MuI._1719_ ),
    .X(\MuI._1734_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5902_  (.A(\MuI._1733_ ),
    .B(\MuI._1734_ ),
    .Y(\MuI._1735_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5903_  (.A_N(\MuI._1698_ ),
    .B(\MuI._1700_ ),
    .X(\MuI._1737_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._5904_  (.A1(\MuI._0750_ ),
    .A2(\MuI._1685_ ),
    .A3(\MuI._1686_ ),
    .B1(\MuI._1696_ ),
    .X(\MuI._1738_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5905_  (.A(\MuI._0755_ ),
    .B(\MuI._0756_ ),
    .Y(\MuI._1739_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5906_  (.A(\MuI._1738_ ),
    .B(\MuI._1739_ ),
    .Y(\MuI._1740_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5907_  (.A(\MuI._1673_ ),
    .B(\MuI._1674_ ),
    .X(\MuI._1741_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5908_  (.A(\MuI._1675_ ),
    .B(\MuI._1677_ ),
    .X(\MuI._1742_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5909_  (.A(\MuI._0685_ ),
    .B(\MuI._1690_ ),
    .C(\MuI._1691_ ),
    .X(\MuI._1743_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5910_  (.A(\MuI._1689_ ),
    .B_N(\MuI._1694_ ),
    .X(\MuI._1744_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5911_  (.A(\MuI._0701_ ),
    .B(\MuI._0704_ ),
    .Y(\MuI._1745_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5912_  (.A1(\MuI._1743_ ),
    .A2(\MuI._1744_ ),
    .B1(\MuI._1745_ ),
    .X(\MuI._1746_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5913_  (.A(\MuI._1743_ ),
    .B(\MuI._1744_ ),
    .C(\MuI._1745_ ),
    .Y(\MuI._1748_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5914_  (.A1(\MuI._1741_ ),
    .A2(\MuI._1742_ ),
    .B1(\MuI._1746_ ),
    .C1(\MuI._1748_ ),
    .X(\MuI._1749_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5915_  (.A1(\MuI._1746_ ),
    .A2(\MuI._1748_ ),
    .B1(\MuI._1741_ ),
    .C1(\MuI._1742_ ),
    .X(\MuI._1750_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5916_  (.A(\MuI._1749_ ),
    .B_N(\MuI._1750_ ),
    .X(\MuI._1751_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5917_  (.A(\MuI._1740_ ),
    .B(\MuI._1751_ ),
    .Y(\MuI._1752_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5918_  (.A(\MuI._1737_ ),
    .B(\MuI._1752_ ),
    .Y(\MuI._1753_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5919_  (.A(\MuI._1735_ ),
    .B(\MuI._1753_ ),
    .X(\MuI._1754_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5920_  (.A(\MuI._1717_ ),
    .B(\MuI._1754_ ),
    .Y(\MuI._1755_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5921_  (.A(\MuI._1716_ ),
    .B(\MuI._1755_ ),
    .Y(\MuI._1756_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._5922_  (.A1(\MuI._1649_ ),
    .A2(\MuI._1708_ ),
    .B1_N(\MuI._1707_ ),
    .Y(\MuI._1757_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5923_  (.A(\MuI._1756_ ),
    .B(\MuI._1757_ ),
    .Y(\MuI._1759_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5924_  (.A(\MuI._1713_ ),
    .B(\MuI._1759_ ),
    .Y(\MuI._1760_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5925_  (.A(\MuI._1712_ ),
    .B(\MuI._1760_ ),
    .X(\MuI._1761_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5926_  (.A(\MuI._1646_ ),
    .B(\MuI._1711_ ),
    .X(\MuI._1762_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5927_  (.A1(\MuI._1713_ ),
    .A2(\MuI._1762_ ),
    .B1(\MuI._1759_ ),
    .X(\MuI._1763_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5928_  (.A1(\MuI._1556_ ),
    .A2(\MuI._1643_ ),
    .B1(\MuI._1641_ ),
    .X(\MuI._1764_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5929_  (.A(\MuI._1761_ ),
    .B(\MuI._1764_ ),
    .X(\MuI._1765_ ));
 sky130_fd_sc_hd__o311a_1 \MuI._5930_  (.A1(\MuI._1460_ ),
    .A2(\MuI._1645_ ),
    .A3(\MuI._1761_ ),
    .B1(\MuI._1763_ ),
    .C1(\MuI._1765_ ),
    .X(\MuI._1766_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._5931_  (.A(\MuI._1717_ ),
    .B_N(\MuI._1754_ ),
    .X(\MuI._1767_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5932_  (.A1(\MuI._1716_ ),
    .A2(\MuI._1755_ ),
    .B1_N(\MuI._1767_ ),
    .X(\MuI._1768_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5933_  (.A(\MuI._1731_ ),
    .B(\MuI._1733_ ),
    .Y(\MuI._1770_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5934_  (.A(\MuI._1737_ ),
    .B(\MuI._1752_ ),
    .Y(\MuI._1771_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5935_  (.A(\MuI._1735_ ),
    .B(\MuI._1753_ ),
    .Y(\MuI._1772_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5936_  (.A(\MuI._1724_ ),
    .Y(\MuI._1773_ ));
 sky130_fd_sc_hd__or4_1 \MuI._5937_  (.A(\MuI._0727_ ),
    .B(\MuI._1724_ ),
    .C(\MuI._1726_ ),
    .D(\MuI._1728_ ),
    .X(\MuI._1774_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5938_  (.A1(\MuI._1743_ ),
    .A2(\MuI._1744_ ),
    .B1(\MuI._1745_ ),
    .Y(\MuI._1775_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5939_  (.A1(\MuI._0725_ ),
    .A2(\MuI._0726_ ),
    .B1(\MuI._0732_ ),
    .Y(\MuI._1776_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5940_  (.A1(\MuI._1775_ ),
    .A2(\MuI._1749_ ),
    .B1(\MuI._1776_ ),
    .C1(\MuI._0733_ ),
    .X(\MuI._1777_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5941_  (.A1(\MuI._0733_ ),
    .A2(\MuI._1776_ ),
    .B1(\MuI._1749_ ),
    .C1(\MuI._1775_ ),
    .Y(\MuI._1778_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5942_  (.A1(\MuI._1773_ ),
    .A2(\MuI._1774_ ),
    .B1(\MuI._1777_ ),
    .C1(\MuI._1778_ ),
    .Y(\MuI._1779_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5943_  (.A1(\MuI._1777_ ),
    .A2(\MuI._1778_ ),
    .B1(\MuI._1773_ ),
    .C1(\MuI._1774_ ),
    .X(\MuI._1781_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5944_  (.A(\MuI._1779_ ),
    .B(\MuI._1781_ ),
    .X(\MuI._1782_ ));
 sky130_fd_sc_hd__a2bb2oi_1 \MuI._5945_  (.A1_N(\MuI._0760_ ),
    .A2_N(\MuI._0761_ ),
    .B1(\MuI._0707_ ),
    .B2(\MuI._0762_ ),
    .Y(\MuI._1783_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5946_  (.A(\MuI._1740_ ),
    .B(\MuI._1751_ ),
    .X(\MuI._1784_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5947_  (.A(\MuI._1738_ ),
    .B(\MuI._1739_ ),
    .Y(\MuI._1785_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5948_  (.A1(\MuI._0763_ ),
    .A2(\MuI._1783_ ),
    .B1(\MuI._1784_ ),
    .C1(\MuI._1785_ ),
    .Y(\MuI._1786_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5949_  (.A1(\MuI._1785_ ),
    .A2(\MuI._1784_ ),
    .B1(\MuI._1783_ ),
    .C1(\MuI._0763_ ),
    .X(\MuI._1787_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._5950_  (.A_N(\MuI._1782_ ),
    .B(\MuI._1786_ ),
    .C(\MuI._1787_ ),
    .Y(\MuI._1788_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5951_  (.A1(\MuI._1787_ ),
    .A2(\MuI._1786_ ),
    .B1_N(\MuI._1782_ ),
    .X(\MuI._1789_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._5952_  (.A1(\MuI._1771_ ),
    .A2(\MuI._1772_ ),
    .B1(\MuI._1788_ ),
    .C1(\MuI._1789_ ),
    .X(\MuI._1790_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._5953_  (.A1(\MuI._1788_ ),
    .A2(\MuI._1789_ ),
    .B1(\MuI._1771_ ),
    .C1(\MuI._1772_ ),
    .Y(\MuI._1792_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5954_  (.A(\MuI._1790_ ),
    .B(\MuI._1792_ ),
    .Y(\MuI._1793_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5955_  (.A(\MuI._1770_ ),
    .B(\MuI._1793_ ),
    .X(\MuI._1794_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5956_  (.A(\MuI._1768_ ),
    .B(\MuI._1794_ ),
    .Y(\MuI._1795_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._5957_  (.A1(\MuI._1777_ ),
    .A2(\MuI._1779_ ),
    .B1(\MuI._0730_ ),
    .Y(\MuI._1796_ ));
 sky130_fd_sc_hd__or3_1 \MuI._5958_  (.A(\MuI._0730_ ),
    .B(\MuI._1777_ ),
    .C(\MuI._1779_ ),
    .X(\MuI._1797_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5959_  (.A(\MuI._1796_ ),
    .B(\MuI._1797_ ),
    .X(\MuI._1798_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5960_  (.A_N(\MuI._0765_ ),
    .B(\MuI._0766_ ),
    .X(\MuI._1799_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5961_  (.A1(\MuI._0737_ ),
    .A2(\MuI._0767_ ),
    .B1(\MuI._1799_ ),
    .Y(\MuI._1800_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5962_  (.A1(\MuI._1787_ ),
    .A2(\MuI._1788_ ),
    .B1(\MuI._1800_ ),
    .C1(\MuI._0769_ ),
    .X(\MuI._1801_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._5963_  (.A1(\MuI._0769_ ),
    .A2(\MuI._1800_ ),
    .B1(\MuI._1788_ ),
    .C1(\MuI._1787_ ),
    .Y(\MuI._1803_ ));
 sky130_fd_sc_hd__and3_1 \MuI._5964_  (.A(\MuI._1798_ ),
    .B(\MuI._1801_ ),
    .C(\MuI._1803_ ),
    .X(\MuI._1804_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._5965_  (.A1(\MuI._1801_ ),
    .A2(\MuI._1803_ ),
    .B1(\MuI._1798_ ),
    .Y(\MuI._1805_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5966_  (.A(\MuI._1804_ ),
    .B(\MuI._1805_ ),
    .Y(\MuI._1806_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5967_  (.A1(\MuI._1770_ ),
    .A2(\MuI._1793_ ),
    .B1(\MuI._1790_ ),
    .X(\MuI._1807_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5968_  (.A(\MuI._1806_ ),
    .B(\MuI._1807_ ),
    .Y(\MuI._1808_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._5969_  (.A(\MuI._1795_ ),
    .B(\MuI._1808_ ),
    .X(\MuI._1809_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5970_  (.A(\MuI._1768_ ),
    .B(\MuI._1794_ ),
    .X(\MuI._1810_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5971_  (.A(\MuI._1756_ ),
    .B(\MuI._1757_ ),
    .Y(\MuI._1811_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5972_  (.A1(\MuI._1795_ ),
    .A2(\MuI._1810_ ),
    .B1(\MuI._1811_ ),
    .X(\MuI._1812_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5973_  (.A(\MuI._1811_ ),
    .B(\MuI._1795_ ),
    .C(\MuI._1810_ ),
    .Y(\MuI._1814_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5974_  (.A(\MuI._1812_ ),
    .B(\MuI._1814_ ),
    .X(\MuI._1815_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5975_  (.A(\MuI._1809_ ),
    .B(\MuI._1815_ ),
    .Y(\MuI._1816_ ));
 sky130_fd_sc_hd__xnor2_4 \MuI._5976_  (.A(\MuI._0740_ ),
    .B(\MuI._0778_ ),
    .Y(\MuI._1817_ ));
 sky130_fd_sc_hd__inv_2 \MuI._5977_  (.A(\MuI._1796_ ),
    .Y(\MuI._1818_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._5978_  (.A1(\MuI._1798_ ),
    .A2(\MuI._1803_ ),
    .B1_N(\MuI._1801_ ),
    .X(\MuI._1819_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5979_  (.A1(\MuI._0771_ ),
    .A2(\MuI._0772_ ),
    .B1(\MuI._0774_ ),
    .X(\MuI._1820_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5980_  (.A(\MuI._0775_ ),
    .B(\MuI._1820_ ),
    .X(\MuI._1821_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._5981_  (.A(\MuI._1819_ ),
    .B(\MuI._1821_ ),
    .X(\MuI._1822_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5982_  (.A(\MuI._1819_ ),
    .B(\MuI._1821_ ),
    .X(\MuI._1823_ ));
 sky130_fd_sc_hd__a21oi_4 \MuI._5983_  (.A1(\MuI._1818_ ),
    .A2(\MuI._1822_ ),
    .B1(\MuI._1823_ ),
    .Y(\MuI._1825_ ));
 sky130_fd_sc_hd__xnor2_4 \MuI._5984_  (.A(\MuI._1817_ ),
    .B(\MuI._1825_ ),
    .Y(\MuI._1826_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._5985_  (.A(\MuI._1806_ ),
    .B(\MuI._1807_ ),
    .Y(\MuI._1827_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5986_  (.A(\MuI._1818_ ),
    .B(\MuI._1822_ ),
    .Y(\MuI._1828_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._5987_  (.A(\MuI._1827_ ),
    .B(\MuI._1828_ ),
    .Y(\MuI._1829_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5988_  (.A(\MuI._1826_ ),
    .B(\MuI._1829_ ),
    .X(\MuI._1830_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._5989_  (.A1(\MuI._1795_ ),
    .A2(\MuI._1814_ ),
    .B1(\MuI._1808_ ),
    .X(\MuI._1831_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._5990_  (.A1(\MuI._1817_ ),
    .A2(\MuI._1825_ ),
    .B1(\MuI._1828_ ),
    .C1(\MuI._1827_ ),
    .X(\MuI._1832_ ));
 sky130_fd_sc_hd__or2_1 \MuI._5991_  (.A(\MuI._1817_ ),
    .B(\MuI._1825_ ),
    .X(\MuI._1833_ ));
 sky130_fd_sc_hd__o311a_1 \MuI._5992_  (.A1(\MuI._1826_ ),
    .A2(\MuI._1829_ ),
    .A3(\MuI._1831_ ),
    .B1(\MuI._1832_ ),
    .C1(\MuI._1833_ ),
    .X(\MuI._1834_ ));
 sky130_fd_sc_hd__o31a_2 \MuI._5993_  (.A1(\MuI._1766_ ),
    .A2(\MuI._1816_ ),
    .A3(\MuI._1830_ ),
    .B1(\MuI._1834_ ),
    .X(\MuI._1836_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._5994_  (.A_N(\MuI._0672_ ),
    .B(\MuI._0783_ ),
    .X(\MuI._1837_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5995_  (.A(\MuI._0673_ ),
    .B(\MuI._0781_ ),
    .X(\MuI._1838_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._5996_  (.A(\MuI._0782_ ),
    .B(\MuI._1838_ ),
    .Y(\MuI._1839_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._5997_  (.A(\MuI._0551_ ),
    .B(\MuI._1837_ ),
    .C(\MuI._1839_ ),
    .Y(\MuI._1840_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._5998_  (.A(\MuI._1836_ ),
    .B(\MuI._1840_ ),
    .C_N(\MuI._0283_ ),
    .X(\MuI._1841_ ));
 sky130_fd_sc_hd__and2_1 \MuI._5999_  (.A(\MuI._3037_ ),
    .B(\MuI._3156_ ),
    .X(\MuI._1842_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6000_  (.A(\MuI._3121_ ),
    .B(\MuI._3123_ ),
    .Y(\MuI._1843_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6001_  (.A_N(\MuI._3110_ ),
    .B(\MuI._3109_ ),
    .X(\MuI._1844_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6002_  (.A1(\MuI._3111_ ),
    .A2(\MuI._3117_ ),
    .B1(\MuI._1844_ ),
    .Y(\MuI._1845_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6003_  (.A(\MuI._1843_ ),
    .B(\MuI._1845_ ),
    .X(\MuI._1847_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6004_  (.A1(\MuI._3113_ ),
    .A2(\MuI._3116_ ),
    .B1_N(\MuI._3114_ ),
    .X(\MuI._1848_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6005_  (.A(\MuI._1847_ ),
    .B(\MuI._1848_ ),
    .X(\MuI._1849_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6006_  (.A(\MuI._3142_ ),
    .B(\MuI._3145_ ),
    .Y(\MuI._1850_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6007_  (.A(\MuI._3094_ ),
    .B(\MuI._3096_ ),
    .Y(\MuI._1851_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6008_  (.A1(\MuI._3135_ ),
    .A2(\MuI._3137_ ),
    .B1_N(\MuI._3136_ ),
    .X(\MuI._1852_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6009_  (.A(\MuI._1274_ ),
    .B(\MuI._2849_ ),
    .Y(\MuI._1853_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6010_  (.A(\MuI._2550_ ),
    .B(\MuI._2517_ ),
    .C(\MuI._2066_ ),
    .D(\MuI._2916_ ),
    .X(\MuI._1854_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6011_  (.A1(\MuI._1813_ ),
    .A2(\MuI._2066_ ),
    .B1(\MuI._2916_ ),
    .B2(\MuI._1318_ ),
    .Y(\MuI._1855_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6012_  (.A(\MuI._1854_ ),
    .B(\MuI._1855_ ),
    .Y(\MuI._1856_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6013_  (.A(\MuI._1853_ ),
    .B(\MuI._1856_ ),
    .Y(\MuI._1858_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6014_  (.A(\MuI._1852_ ),
    .B(\MuI._1858_ ),
    .Y(\MuI._1859_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6015_  (.A(\MuI._1851_ ),
    .B(\MuI._1859_ ),
    .Y(\MuI._1860_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6016_  (.A(\MuI._3098_ ),
    .B(\MuI._3100_ ),
    .X(\MuI._1861_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6017_  (.A(\MuI._1860_ ),
    .B(\MuI._1861_ ),
    .X(\MuI._1862_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6018_  (.A(\MuI._0878_ ),
    .B(\MuI._2789_ ),
    .C(\MuI._3107_ ),
    .X(\MuI._1863_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6019_  (.A(\MuI._0878_ ),
    .B(\MuI._2797_ ),
    .Y(\MuI._1864_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6020_  (.A(\MuI._0735_ ),
    .B(\MuI._1153_ ),
    .C(\MuI._2682_ ),
    .D(\MuI._2594_ ),
    .X(\MuI._1865_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6021_  (.A1(\MuI._1153_ ),
    .A2(\MuI._2914_ ),
    .B1(\MuI._2594_ ),
    .B2(\MuI._0746_ ),
    .Y(\MuI._1866_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6022_  (.A(\MuI._1865_ ),
    .B(\MuI._1866_ ),
    .Y(\MuI._1867_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6023_  (.A(\MuI._1864_ ),
    .B(\MuI._1867_ ),
    .Y(\MuI._1869_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6024_  (.A1(\MuI._3105_ ),
    .A2(\MuI._1863_ ),
    .B1(\MuI._1869_ ),
    .X(\MuI._1870_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6025_  (.A(\MuI._3105_ ),
    .B(\MuI._1863_ ),
    .C(\MuI._1869_ ),
    .Y(\MuI._1871_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6026_  (.A(\MuI._1870_ ),
    .B(\MuI._1871_ ),
    .Y(\MuI._1872_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6027_  (.A1(\MuI._0625_ ),
    .A2(\MuI._2789_ ),
    .B1(\MuI._2791_ ),
    .B2(\MuI._0372_ ),
    .Y(\MuI._1873_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6028_  (.A(\MuI._0372_ ),
    .B(\MuI._0614_ ),
    .C(\MuI._2789_ ),
    .D(\MuI._2791_ ),
    .X(\MuI._1874_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6029_  (.A(\MuI._1873_ ),
    .B(\MuI._1874_ ),
    .Y(\MuI._1875_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6030_  (.A(\MuI._2787_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._1876_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6031_  (.A(\MuI._1875_ ),
    .B(\MuI._1876_ ),
    .Y(\MuI._1877_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6032_  (.A(\MuI._1872_ ),
    .B(\MuI._1877_ ),
    .Y(\MuI._1878_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6033_  (.A(\MuI._1862_ ),
    .B(\MuI._1878_ ),
    .Y(\MuI._1880_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6034_  (.A(\MuI._1850_ ),
    .B(\MuI._1880_ ),
    .X(\MuI._1881_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6035_  (.A(\MuI._3103_ ),
    .B_N(\MuI._3119_ ),
    .X(\MuI._1882_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6036_  (.A(\MuI._1881_ ),
    .B(\MuI._1882_ ),
    .Y(\MuI._1883_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6037_  (.A(\MuI._3133_ ),
    .B(\MuI._3140_ ),
    .Y(\MuI._1884_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6038_  (.A(\MuI._1884_ ),
    .Y(\MuI._1885_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6039_  (.A(\MuI._0581_ ),
    .B(\MuI._2851_ ),
    .Y(\MuI._1886_ ));
 sky130_fd_sc_hd__and2_2 \MuI._6040_  (.A(\MuI._0339_ ),
    .B(\MuI._2975_ ),
    .X(\MuI._1887_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6041_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._2976_ ),
    .X(\MuI._1888_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6042_  (.A(\MuI._1887_ ),
    .B(\MuI._1888_ ),
    .X(\MuI._1889_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6043_  (.A(\MuI._1886_ ),
    .B(\MuI._1889_ ),
    .Y(\MuI._1891_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6044_  (.A(\MuI._3129_ ),
    .B(\MuI._3131_ ),
    .Y(\MuI._1892_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6045_  (.A(\MuI._1891_ ),
    .B(\MuI._1892_ ),
    .X(\MuI._1893_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6046_  (.A(\MuI._1483_ ),
    .B(\MuI._2583_ ),
    .Y(\MuI._1894_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6047_  (.A(\MuI._0779_ ),
    .B(\MuI._1021_ ),
    .C(\MuI._2704_ ),
    .D(\MuI._2649_ ),
    .X(\MuI._1895_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6048_  (.A1(\MuI._1032_ ),
    .A2(\MuI._2800_ ),
    .B1(\MuI._2919_ ),
    .B2(\MuI._0790_ ),
    .Y(\MuI._1896_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6049_  (.A(\MuI._1895_ ),
    .B(\MuI._1896_ ),
    .Y(\MuI._1897_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6050_  (.A(\MuI._1894_ ),
    .B(\MuI._1897_ ),
    .Y(\MuI._1898_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6051_  (.A(\MuI._1893_ ),
    .B(\MuI._1898_ ),
    .X(\MuI._1899_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6052_  (.A(\MuI._3067_ ),
    .B(\MuI._1899_ ),
    .Y(\MuI._1900_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6053_  (.A(\MuI._1885_ ),
    .B(\MuI._1900_ ),
    .Y(\MuI._1902_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6054_  (.A(\MuI._3147_ ),
    .B(\MuI._1902_ ),
    .X(\MuI._1903_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6055_  (.A(\MuI._1883_ ),
    .B(\MuI._1903_ ),
    .X(\MuI._1904_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6056_  (.A(\MuI._3149_ ),
    .B(\MuI._3151_ ),
    .Y(\MuI._1905_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6057_  (.A1(\MuI._3125_ ),
    .A2(\MuI._3152_ ),
    .B1(\MuI._1905_ ),
    .X(\MuI._1906_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6058_  (.A(\MuI._1904_ ),
    .B(\MuI._1906_ ),
    .Y(\MuI._1907_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._6059_  (.A(\MuI._1849_ ),
    .B(\MuI._1907_ ),
    .Y(\MuI._1908_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6060_  (.A1(\MuI._3154_ ),
    .A2(\MuI._1842_ ),
    .B1(\MuI._1908_ ),
    .Y(\MuI._1909_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6061_  (.A_N(\MuI._3036_ ),
    .B(\MuI._3035_ ),
    .X(\MuI._1910_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6062_  (.A(\MuI._3033_ ),
    .B(\MuI._1910_ ),
    .Y(\MuI._1911_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6063_  (.A(\MuI._3154_ ),
    .B(\MuI._1842_ ),
    .C(\MuI._1908_ ),
    .X(\MuI._1913_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6064_  (.A(\MuI._1909_ ),
    .B(\MuI._1913_ ),
    .X(\MuI._1914_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6065_  (.A(\MuI._1911_ ),
    .B_N(\MuI._1914_ ),
    .X(\MuI._1915_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6066_  (.A(\MuI._1848_ ),
    .B_N(\MuI._1847_ ),
    .X(\MuI._1916_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._6067_  (.A1(\MuI._1843_ ),
    .A2(\MuI._1845_ ),
    .B1(\MuI._1916_ ),
    .Y(\MuI._1917_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6068_  (.A(\MuI._1850_ ),
    .B(\MuI._1880_ ),
    .X(\MuI._1918_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6069_  (.A1(\MuI._1881_ ),
    .A2(\MuI._1882_ ),
    .B1(\MuI._1918_ ),
    .Y(\MuI._1919_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6070_  (.A1(\MuI._1872_ ),
    .A2(\MuI._1877_ ),
    .B1(\MuI._1870_ ),
    .Y(\MuI._1920_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6071_  (.A(\MuI._1919_ ),
    .B(\MuI._1920_ ),
    .X(\MuI._1921_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6072_  (.A1(\MuI._1873_ ),
    .A2(\MuI._1876_ ),
    .B1_N(\MuI._1874_ ),
    .X(\MuI._1922_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6073_  (.A(\MuI._1921_ ),
    .B(\MuI._1922_ ),
    .Y(\MuI._1924_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6074_  (.A(\MuI._3067_ ),
    .B(\MuI._1899_ ),
    .Y(\MuI._1925_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6075_  (.A1(\MuI._1885_ ),
    .A2(\MuI._1900_ ),
    .B1(\MuI._1925_ ),
    .Y(\MuI._1926_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6076_  (.A(\MuI._1852_ ),
    .B_N(\MuI._1858_ ),
    .X(\MuI._1927_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6077_  (.A(\MuI._1851_ ),
    .B(\MuI._1859_ ),
    .Y(\MuI._1928_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6078_  (.A1(\MuI._1285_ ),
    .A2(\MuI._2849_ ),
    .A3(\MuI._1856_ ),
    .B1(\MuI._1854_ ),
    .X(\MuI._1929_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6079_  (.A1(\MuI._1894_ ),
    .A2(\MuI._1896_ ),
    .B1_N(\MuI._1895_ ),
    .X(\MuI._1930_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6080_  (.A(\MuI._2473_ ),
    .B(\MuI._3091_ ),
    .Y(\MuI._1931_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6081_  (.A(\MuI._1472_ ),
    .B(\MuI._1296_ ),
    .C(\MuI._1791_ ),
    .D(\MuI._2055_ ),
    .X(\MuI._1932_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6082_  (.A1(\MuI._1472_ ),
    .A2(\MuI._1802_ ),
    .B1(\MuI._2843_ ),
    .B2(\MuI._1307_ ),
    .Y(\MuI._1933_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6083_  (.A(\MuI._1932_ ),
    .B(\MuI._1933_ ),
    .Y(\MuI._1935_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6084_  (.A(\MuI._1931_ ),
    .B(\MuI._1935_ ),
    .Y(\MuI._1936_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6085_  (.A(\MuI._1930_ ),
    .B(\MuI._1936_ ),
    .Y(\MuI._1937_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6086_  (.A(\MuI._1929_ ),
    .B(\MuI._1937_ ),
    .Y(\MuI._1938_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6087_  (.A1(\MuI._1927_ ),
    .A2(\MuI._1928_ ),
    .B1(\MuI._1938_ ),
    .X(\MuI._1939_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6088_  (.A(\MuI._1927_ ),
    .B(\MuI._1928_ ),
    .C(\MuI._1938_ ),
    .Y(\MuI._1940_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6089_  (.A(\MuI._1939_ ),
    .B(\MuI._1940_ ),
    .Y(\MuI._1941_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6090_  (.A(\MuI._0867_ ),
    .B(\MuI._2594_ ),
    .Y(\MuI._1942_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6091_  (.A(\MuI._0735_ ),
    .B(\MuI._2813_ ),
    .C(\MuI._2627_ ),
    .D(\MuI._2682_ ),
    .X(\MuI._1943_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6092_  (.A1(\MuI._1153_ ),
    .A2(\MuI._2627_ ),
    .B1(\MuI._2914_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._1944_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6093_  (.A(\MuI._1943_ ),
    .B(\MuI._1944_ ),
    .Y(\MuI._1946_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6094_  (.A(\MuI._1942_ ),
    .B(\MuI._1946_ ),
    .Y(\MuI._1947_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6095_  (.A1(\MuI._1864_ ),
    .A2(\MuI._1866_ ),
    .B1_N(\MuI._1865_ ),
    .X(\MuI._1948_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6096_  (.A(\MuI._1947_ ),
    .B(\MuI._1948_ ),
    .Y(\MuI._1949_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6097_  (.A1(\MuI._0625_ ),
    .A2(\MuI._2797_ ),
    .B1(\MuI._2789_ ),
    .B2(\MuI._0372_ ),
    .Y(\MuI._1950_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6098_  (.A(\MuI._0372_ ),
    .B(\MuI._0625_ ),
    .C(\MuI._2797_ ),
    .D(\MuI._2789_ ),
    .X(\MuI._1951_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6099_  (.A(\MuI._1950_ ),
    .B(\MuI._1951_ ),
    .Y(\MuI._1952_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6100_  (.A(\MuI._2791_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._1953_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6101_  (.A(\MuI._1952_ ),
    .B(\MuI._1953_ ),
    .Y(\MuI._1954_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6102_  (.A(\MuI._1949_ ),
    .B(\MuI._1954_ ),
    .Y(\MuI._1955_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6103_  (.A(\MuI._1941_ ),
    .B(\MuI._1955_ ),
    .Y(\MuI._1957_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6104_  (.A(\MuI._1926_ ),
    .B(\MuI._1957_ ),
    .Y(\MuI._1958_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6105_  (.A(\MuI._1860_ ),
    .B(\MuI._1861_ ),
    .X(\MuI._1959_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6106_  (.A(\MuI._1860_ ),
    .B(\MuI._1861_ ),
    .Y(\MuI._1960_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6107_  (.A1(\MuI._1959_ ),
    .A2(\MuI._1878_ ),
    .B1_N(\MuI._1960_ ),
    .Y(\MuI._1961_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6108_  (.A(\MuI._1958_ ),
    .B(\MuI._1961_ ),
    .Y(\MuI._1962_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6109_  (.A(\MuI._1891_ ),
    .B(\MuI._1892_ ),
    .Y(\MuI._1963_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6110_  (.A(\MuI._1893_ ),
    .B(\MuI._1898_ ),
    .Y(\MuI._1964_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6111_  (.A1(\MuI._0339_ ),
    .A2(\MuI._2851_ ),
    .B1(\MuI._2975_ ),
    .B2(\MuI._0515_ ),
    .Y(\MuI._1965_ ));
 sky130_fd_sc_hd__a31oi_2 \MuI._6112_  (.A1(\MuI._2851_ ),
    .A2(\MuI._0526_ ),
    .A3(\MuI._1887_ ),
    .B1(\MuI._1965_ ),
    .Y(\MuI._1966_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6113_  (.A(\MuI._1887_ ),
    .B(\MuI._1888_ ),
    .X(\MuI._1968_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6114_  (.A1(\MuI._0581_ ),
    .A2(\MuI._2851_ ),
    .A3(\MuI._1889_ ),
    .B1(\MuI._1968_ ),
    .X(\MuI._1969_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6115_  (.A(\MuI._1966_ ),
    .B(\MuI._1969_ ),
    .X(\MuI._1970_ ));
 sky130_fd_sc_hd__nand2_2 \MuI._6116_  (.A(\MuI._1021_ ),
    .B(\MuI.b_operand[14] ),
    .Y(\MuI._1971_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6117_  (.A(\MuI._0559_ ),
    .B(\MuI._0768_ ),
    .C(\MuI._2693_ ),
    .D(\MuI._2638_ ),
    .X(\MuI._1972_ ));
 sky130_fd_sc_hd__a22oi_2 \MuI._6118_  (.A1(\MuI._0779_ ),
    .A2(\MuI._2802_ ),
    .B1(\MuI._2803_ ),
    .B2(\MuI._2894_ ),
    .Y(\MuI._1973_ ));
 sky130_fd_sc_hd__nor2_2 \MuI._6119_  (.A(\MuI._1972_ ),
    .B(\MuI._1973_ ),
    .Y(\MuI._1974_ ));
 sky130_fd_sc_hd__xnor2_4 \MuI._6120_  (.A(\MuI._1971_ ),
    .B(\MuI._1974_ ),
    .Y(\MuI._1975_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6121_  (.A(\MuI._1970_ ),
    .B(\MuI._1975_ ),
    .Y(\MuI._1976_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6122_  (.A1(\MuI._1963_ ),
    .A2(\MuI._1964_ ),
    .B1(\MuI._1976_ ),
    .Y(\MuI._1977_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6123_  (.A(\MuI._1963_ ),
    .B(\MuI._1964_ ),
    .C(\MuI._1976_ ),
    .X(\MuI._1979_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6124_  (.A(\MuI._1977_ ),
    .B(\MuI._1979_ ),
    .Y(\MuI._1980_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6125_  (.A(\MuI._1962_ ),
    .B(\MuI._1980_ ),
    .Y(\MuI._1981_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6126_  (.A(\MuI._1883_ ),
    .B_N(\MuI._1903_ ),
    .X(\MuI._1982_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6127_  (.A1(\MuI._3147_ ),
    .A2(\MuI._1902_ ),
    .B1(\MuI._1982_ ),
    .X(\MuI._1983_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6128_  (.A(\MuI._1981_ ),
    .B(\MuI._1983_ ),
    .Y(\MuI._1984_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6129_  (.A(\MuI._1924_ ),
    .B(\MuI._1984_ ),
    .Y(\MuI._1985_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6130_  (.A(\MuI._1904_ ),
    .B_N(\MuI._1906_ ),
    .X(\MuI._1986_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6131_  (.A(\MuI._1849_ ),
    .B_N(\MuI._1907_ ),
    .X(\MuI._1987_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6132_  (.A(\MuI._1986_ ),
    .B(\MuI._1987_ ),
    .X(\MuI._1988_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6133_  (.A(\MuI._1985_ ),
    .B(\MuI._1988_ ),
    .Y(\MuI._1990_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6134_  (.A(\MuI._1985_ ),
    .B(\MuI._1988_ ),
    .X(\MuI._1991_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6135_  (.A(\MuI._1990_ ),
    .B(\MuI._1991_ ),
    .Y(\MuI._1992_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._6136_  (.A(\MuI._1917_ ),
    .B(\MuI._1992_ ),
    .Y(\MuI._1993_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6137_  (.A1(\MuI._1909_ ),
    .A2(\MuI._1915_ ),
    .B1(\MuI._1993_ ),
    .Y(\MuI._1994_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6138_  (.A(\MuI._1993_ ),
    .B(\MuI._1909_ ),
    .C(\MuI._1915_ ),
    .X(\MuI._1995_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6139_  (.A(\MuI._1994_ ),
    .B(\MuI._1995_ ),
    .Y(\MuI._1996_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6140_  (.A_N(\MuI._3180_ ),
    .B(\MuI._2960_ ),
    .X(\MuI._1997_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6141_  (.A1(\MuI._3157_ ),
    .A2(\MuI._3179_ ),
    .B1_N(\MuI._1997_ ),
    .X(\MuI._1998_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6142_  (.A(\MuI._1911_ ),
    .B(\MuI._1914_ ),
    .Y(\MuI._1999_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6143_  (.A(\MuI._1998_ ),
    .B_N(\MuI._1999_ ),
    .X(\MuI._2001_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6144_  (.A(\MuI._2001_ ),
    .Y(\MuI._2002_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6145_  (.A_N(\MuI._1999_ ),
    .B(\MuI._1998_ ),
    .X(\MuI._2003_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6146_  (.A(\MuI._2002_ ),
    .B(\MuI._2003_ ),
    .Y(\MuI._2004_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6147_  (.A(\MuI._1996_ ),
    .B(\MuI._2004_ ),
    .Y(\MuI._2005_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6148_  (.A(\MuI.a_operand[22] ),
    .B(\MuI._2693_ ),
    .C(\MuI._2638_ ),
    .X(\MuI._2006_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6149_  (.A(\MuI._0504_ ),
    .B(\MuI._2006_ ),
    .X(\MuI._2007_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6150_  (.A(\MuI._0328_ ),
    .B(\MuI._2802_ ),
    .X(\MuI._2008_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6151_  (.A1(\MuI.a_operand[25] ),
    .A2(\MuI._2889_ ),
    .A3(\MuI._2890_ ),
    .B1(\MuI._2649_ ),
    .X(\MuI._2009_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6152_  (.A1(\MuI._0482_ ),
    .A2(\MuI._0493_ ),
    .B1_N(\MuI._2006_ ),
    .X(\MuI._2010_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._6153_  (.A1(\MuI._2008_ ),
    .A2(\MuI._2009_ ),
    .B1(\MuI._2010_ ),
    .C1(\MuI._0570_ ),
    .D1(\MuI._2583_ ),
    .X(\MuI._2012_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6154_  (.A(\MuI._1032_ ),
    .B(\MuI._2473_ ),
    .Y(\MuI._2013_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6155_  (.A(\MuI._0559_ ),
    .B(\MuI._0768_ ),
    .C(\MuI._3000_ ),
    .D(\MuI._2754_ ),
    .X(\MuI._2014_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6156_  (.A1(\MuI._0779_ ),
    .A2(\MuI._2550_ ),
    .B1(\MuI._2517_ ),
    .B2(\MuI._2894_ ),
    .Y(\MuI._2015_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6157_  (.A(\MuI._2014_ ),
    .B(\MuI._2015_ ),
    .Y(\MuI._2016_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6158_  (.A(\MuI._2013_ ),
    .B(\MuI._2016_ ),
    .Y(\MuI._2017_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6159_  (.A1(\MuI._2007_ ),
    .A2(\MuI._2012_ ),
    .B1(\MuI._2017_ ),
    .Y(\MuI._2018_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6160_  (.A(\MuI._0779_ ),
    .B(\MuI._1010_ ),
    .C(\MuI._3000_ ),
    .D(\MuI._2754_ ),
    .X(\MuI._2019_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6161_  (.A(\MuI._1483_ ),
    .B(\MuI._1263_ ),
    .Y(\MuI._2020_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6162_  (.A1(\MuI._1021_ ),
    .A2(\MuI._2550_ ),
    .B1(\MuI._2517_ ),
    .B2(\MuI._0779_ ),
    .Y(\MuI._2021_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6163_  (.A(\MuI._2019_ ),
    .B(\MuI._2020_ ),
    .C(\MuI._2021_ ),
    .X(\MuI._2023_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6164_  (.A(\MuI._2019_ ),
    .B_N(\MuI._2023_ ),
    .X(\MuI._2024_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6165_  (.A(\MuI._2007_ ),
    .B(\MuI._2012_ ),
    .C(\MuI._2017_ ),
    .X(\MuI._2025_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6166_  (.A(\MuI._2018_ ),
    .B(\MuI._2024_ ),
    .C(\MuI._2025_ ),
    .Y(\MuI._2026_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6167_  (.A1(\MuI._2018_ ),
    .A2(\MuI._2025_ ),
    .B1(\MuI._2024_ ),
    .X(\MuI._2027_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6168_  (.A(\MuI._0790_ ),
    .B(\MuI._2796_ ),
    .Y(\MuI._2028_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6169_  (.A1(\MuI._0570_ ),
    .A2(\MuI._2800_ ),
    .B1(\MuI._2919_ ),
    .B2(\MuI._0339_ ),
    .Y(\MuI._2029_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6170_  (.A(\MuI._0328_ ),
    .B(\MuI._2894_ ),
    .C(\MuI._2802_ ),
    .D(\MuI._2803_ ),
    .X(\MuI._2030_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6171_  (.A1(\MuI._2028_ ),
    .A2(\MuI._2029_ ),
    .B1_N(\MuI._2030_ ),
    .Y(\MuI._2031_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6172_  (.A1(\MuI._2019_ ),
    .A2(\MuI._2021_ ),
    .B1(\MuI._2020_ ),
    .Y(\MuI._2032_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6173_  (.A(\MuI._2023_ ),
    .B(\MuI._2031_ ),
    .C(\MuI._2032_ ),
    .Y(\MuI._2034_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6174_  (.A(\MuI.a_operand[19] ),
    .B(\MuI._1461_ ),
    .C(\MuI._1296_ ),
    .D(\MuI.b_operand[15] ),
    .X(\MuI._2035_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6175_  (.A(\MuI.b_operand[17] ),
    .B(\MuI._2843_ ),
    .Y(\MuI._2036_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6176_  (.A1(\MuI._1461_ ),
    .A2(\MuI._1296_ ),
    .B1(\MuI._1791_ ),
    .B2(\MuI._1010_ ),
    .Y(\MuI._2037_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6177_  (.A(\MuI._2035_ ),
    .B(\MuI._2036_ ),
    .C(\MuI._2037_ ),
    .X(\MuI._2038_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6178_  (.A(\MuI._2035_ ),
    .B_N(\MuI._2038_ ),
    .X(\MuI._2039_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6179_  (.A1(\MuI._2023_ ),
    .A2(\MuI._2032_ ),
    .B1(\MuI._2031_ ),
    .X(\MuI._2040_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6180_  (.A(\MuI._2034_ ),
    .B(\MuI._2039_ ),
    .C(\MuI._2040_ ),
    .Y(\MuI._2041_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6181_  (.A(\MuI._2034_ ),
    .B(\MuI._2041_ ),
    .Y(\MuI._2042_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6182_  (.A(\MuI._2026_ ),
    .B(\MuI._2027_ ),
    .C(\MuI._2042_ ),
    .X(\MuI._2043_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6183_  (.A1(\MuI._2026_ ),
    .A2(\MuI._2027_ ),
    .B1(\MuI._2042_ ),
    .Y(\MuI._2045_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6184_  (.A(\MuI._2817_ ),
    .B(\MuI._3091_ ),
    .Y(\MuI._2046_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6185_  (.A(\MuI._2939_ ),
    .B(\MuI._1142_ ),
    .C(\MuI._1483_ ),
    .D(\MuI._2066_ ),
    .X(\MuI._2047_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._6186_  (.A1(\MuI._2813_ ),
    .A2(\MuI._1483_ ),
    .B1(\MuI._2066_ ),
    .B2(\MuI._2814_ ),
    .X(\MuI._2048_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6187_  (.A_N(\MuI._2047_ ),
    .B(\MuI._2048_ ),
    .X(\MuI._2049_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6188_  (.A(\MuI._2046_ ),
    .B(\MuI._2049_ ),
    .Y(\MuI._2050_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6189_  (.A(\MuI._2939_ ),
    .B(\MuI._2811_ ),
    .C(\MuI._2843_ ),
    .D(\MuI._2840_ ),
    .X(\MuI._2051_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6190_  (.A1(\MuI._2813_ ),
    .A2(\MuI._2066_ ),
    .B1(\MuI._2916_ ),
    .B2(\MuI._2814_ ),
    .Y(\MuI._2052_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._6191_  (.A_N(\MuI._2051_ ),
    .B_N(\MuI._2052_ ),
    .C(\MuI._0867_ ),
    .D(\MuI._2627_ ),
    .X(\MuI._2053_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6192_  (.A(\MuI._2051_ ),
    .B(\MuI._2053_ ),
    .Y(\MuI._2054_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6193_  (.A(\MuI._2050_ ),
    .B(\MuI._2054_ ),
    .Y(\MuI._2056_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6194_  (.A1(\MuI._0614_ ),
    .A2(\MuI._2849_ ),
    .B1(\MuI._2914_ ),
    .B2(\MuI._0361_ ),
    .Y(\MuI._2057_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6195_  (.A(\MuI._0361_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._2849_ ),
    .D(\MuI._2914_ ),
    .X(\MuI._2058_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6196_  (.A(\MuI._2057_ ),
    .B(\MuI._2058_ ),
    .Y(\MuI._2059_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6197_  (.A(\MuI._2594_ ),
    .B(\MuI._0449_ ),
    .Y(\MuI._2060_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6198_  (.A(\MuI._2059_ ),
    .B(\MuI._2060_ ),
    .Y(\MuI._2061_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6199_  (.A(\MuI._2056_ ),
    .B(\MuI._2061_ ),
    .Y(\MuI._2062_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6200_  (.A(\MuI._2043_ ),
    .B(\MuI._2045_ ),
    .C(\MuI._2062_ ),
    .X(\MuI._2063_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6201_  (.A(\MuI._2030_ ),
    .B(\MuI._2029_ ),
    .Y(\MuI._2064_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._6202_  (.A(\MuI._2028_ ),
    .B(\MuI._2064_ ),
    .Y(\MuI._2065_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6203_  (.A1(\MuI._1887_ ),
    .A2(\MuI._2065_ ),
    .B1(\MuI._2851_ ),
    .C1(\MuI._0526_ ),
    .X(\MuI._2067_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6204_  (.A1(\MuI._2008_ ),
    .A2(\MuI._2009_ ),
    .B1(\MuI._2010_ ),
    .X(\MuI._2068_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6205_  (.A1(\MuI._0592_ ),
    .A2(\MuI._2860_ ),
    .B1(\MuI._2068_ ),
    .Y(\MuI._2069_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6206_  (.A(\MuI._2012_ ),
    .B(\MuI._2069_ ),
    .Y(\MuI._2070_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6207_  (.A(\MuI._2067_ ),
    .B(\MuI._2070_ ),
    .X(\MuI._2071_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6208_  (.A1(\MuI._2043_ ),
    .A2(\MuI._2045_ ),
    .B1(\MuI._2062_ ),
    .Y(\MuI._2072_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6209_  (.A(\MuI._2063_ ),
    .B(\MuI._2071_ ),
    .C(\MuI._2072_ ),
    .Y(\MuI._2073_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6210_  (.A1(\MuI._2063_ ),
    .A2(\MuI._2072_ ),
    .B1(\MuI._2071_ ),
    .X(\MuI._2074_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6211_  (.A1(\MuI._2034_ ),
    .A2(\MuI._2040_ ),
    .B1(\MuI._2039_ ),
    .X(\MuI._2075_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6212_  (.A1(\MuI._1274_ ),
    .A2(\MuI._3091_ ),
    .A3(\MuI._1935_ ),
    .B1(\MuI._1932_ ),
    .X(\MuI._2076_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6213_  (.A1(\MuI._2035_ ),
    .A2(\MuI._2037_ ),
    .B1(\MuI._2036_ ),
    .Y(\MuI._2078_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6214_  (.A1(\MuI._1971_ ),
    .A2(\MuI._1973_ ),
    .B1_N(\MuI._1972_ ),
    .Y(\MuI._2079_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6215_  (.A1(\MuI._2038_ ),
    .A2(\MuI._2078_ ),
    .B1(\MuI._2079_ ),
    .X(\MuI._2080_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6216_  (.A(\MuI._2038_ ),
    .B(\MuI._2079_ ),
    .C(\MuI._2078_ ),
    .Y(\MuI._2081_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6217_  (.A1(\MuI._2076_ ),
    .A2(\MuI._2080_ ),
    .B1_N(\MuI._2081_ ),
    .X(\MuI._2082_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6218_  (.A(\MuI._2041_ ),
    .B(\MuI._2075_ ),
    .C(\MuI._2082_ ),
    .X(\MuI._2083_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6219_  (.A1(\MuI._2041_ ),
    .A2(\MuI._2075_ ),
    .B1(\MuI._2082_ ),
    .Y(\MuI._2084_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._6220_  (.A1_N(\MuI._0867_ ),
    .A2_N(\MuI._2849_ ),
    .B1(\MuI._2051_ ),
    .B2(\MuI._2052_ ),
    .X(\MuI._2085_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6221_  (.A(\MuI._2053_ ),
    .B(\MuI._2085_ ),
    .Y(\MuI._2086_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6222_  (.A(\MuI.b_operand[19] ),
    .B(\MuI._2811_ ),
    .C(\MuI._2840_ ),
    .D(\MuI._2616_ ),
    .X(\MuI._2087_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6223_  (.A1(\MuI._1142_ ),
    .A2(\MuI._2916_ ),
    .B1(\MuI._2627_ ),
    .B2(\MuI._2814_ ),
    .Y(\MuI._2089_ ));
 sky130_fd_sc_hd__and4bb_1 \MuI._6224_  (.A_N(\MuI._2087_ ),
    .B_N(\MuI._2089_ ),
    .C(\MuI.b_operand[20] ),
    .D(\MuI._2682_ ),
    .X(\MuI._2090_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6225_  (.A(\MuI._2087_ ),
    .B(\MuI._2090_ ),
    .Y(\MuI._2091_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6226_  (.A(\MuI._2086_ ),
    .B(\MuI._2091_ ),
    .Y(\MuI._2092_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6227_  (.A1(\MuI._0603_ ),
    .A2(\MuI._2914_ ),
    .B1(\MuI._2594_ ),
    .B2(\MuI._2826_ ),
    .Y(\MuI._2093_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6228_  (.A(\MuI._2826_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._2682_ ),
    .D(\MuI._2594_ ),
    .X(\MuI._2094_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6229_  (.A(\MuI._2093_ ),
    .B(\MuI._2094_ ),
    .Y(\MuI._2095_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6230_  (.A(\MuI._2797_ ),
    .B(\MuI._0438_ ),
    .Y(\MuI._2096_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6231_  (.A(\MuI._2095_ ),
    .B(\MuI._2096_ ),
    .Y(\MuI._2097_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6232_  (.A(\MuI._2092_ ),
    .B(\MuI._2097_ ),
    .Y(\MuI._2098_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6233_  (.A(\MuI._2083_ ),
    .B(\MuI._2084_ ),
    .C(\MuI._2098_ ),
    .X(\MuI._2100_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6234_  (.A(\MuI._2083_ ),
    .B_N(\MuI._2100_ ),
    .X(\MuI._2101_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6235_  (.A(\MuI._2073_ ),
    .B(\MuI._2074_ ),
    .C(\MuI._2101_ ),
    .Y(\MuI._2102_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6236_  (.A1(\MuI._2073_ ),
    .A2(\MuI._2074_ ),
    .B1(\MuI._2101_ ),
    .X(\MuI._2103_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6237_  (.A(\MuI._2860_ ),
    .B(\MuI._0515_ ),
    .C(\MuI._2008_ ),
    .X(\MuI._2104_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6238_  (.A1(\MuI._0350_ ),
    .A2(\MuI._2860_ ),
    .B1(\MuI._2800_ ),
    .B2(\MuI._0537_ ),
    .Y(\MuI._2105_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6239_  (.A(\MuI._2104_ ),
    .B(\MuI._2105_ ),
    .Y(\MuI._2106_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6240_  (.A(\MuI._2102_ ),
    .B(\MuI._2103_ ),
    .C(\MuI._2106_ ),
    .Y(\MuI._2107_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6241_  (.A(\MuI._2860_ ),
    .B(\MuI._0537_ ),
    .Y(\MuI._2108_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6242_  (.A(\MuI._2814_ ),
    .B(\MuI._2813_ ),
    .C(\MuI._1021_ ),
    .D(\MuI._1483_ ),
    .X(\MuI._2109_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6243_  (.A1(\MuI._1153_ ),
    .A2(\MuI._1032_ ),
    .B1(\MuI._1483_ ),
    .B2(\MuI._0735_ ),
    .Y(\MuI._2111_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6244_  (.A(\MuI._2109_ ),
    .B(\MuI._2111_ ),
    .Y(\MuI._2112_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6245_  (.A(\MuI._0878_ ),
    .B(\MuI._2077_ ),
    .C(\MuI._2112_ ),
    .X(\MuI._2113_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6246_  (.A1(\MuI._0878_ ),
    .A2(\MuI._2077_ ),
    .B1(\MuI._2112_ ),
    .Y(\MuI._2114_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6247_  (.A(\MuI._2113_ ),
    .B(\MuI._2114_ ),
    .Y(\MuI._2115_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6248_  (.A1(\MuI._0878_ ),
    .A2(\MuI._3091_ ),
    .A3(\MuI._2048_ ),
    .B1(\MuI._2047_ ),
    .X(\MuI._2116_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6249_  (.A(\MuI._2115_ ),
    .B(\MuI._2116_ ),
    .X(\MuI._2117_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6250_  (.A(\MuI._2115_ ),
    .B(\MuI._2116_ ),
    .Y(\MuI._2118_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6251_  (.A(\MuI._2117_ ),
    .B(\MuI._2118_ ),
    .Y(\MuI._2119_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6252_  (.A(\MuI._0361_ ),
    .B(\MuI._0614_ ),
    .C(\MuI._3091_ ),
    .X(\MuI._2120_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._6253_  (.A1(\MuI._0614_ ),
    .A2(\MuI._3091_ ),
    .B1(\MuI._2849_ ),
    .B2(\MuI._0372_ ),
    .X(\MuI._2122_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6254_  (.A1(\MuI._2849_ ),
    .A2(\MuI._2120_ ),
    .B1_N(\MuI._2122_ ),
    .X(\MuI._2123_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6255_  (.A(\MuI._2914_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._2124_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6256_  (.A(\MuI._2123_ ),
    .B(\MuI._2124_ ),
    .X(\MuI._2125_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6257_  (.A(\MuI._2119_ ),
    .B(\MuI._2125_ ),
    .Y(\MuI._2126_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6258_  (.A(\MuI._0790_ ),
    .B(\MuI._1274_ ),
    .Y(\MuI._2127_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6259_  (.A(\MuI._0328_ ),
    .B(\MuI._2894_ ),
    .C(\MuI._2550_ ),
    .D(\MuI._2517_ ),
    .X(\MuI._2128_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6260_  (.A1(\MuI._0570_ ),
    .A2(\MuI._1318_ ),
    .B1(\MuI._1813_ ),
    .B2(\MuI._0339_ ),
    .Y(\MuI._2129_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6261_  (.A(\MuI._2128_ ),
    .B(\MuI._2129_ ),
    .Y(\MuI._2130_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._6262_  (.A(\MuI._2127_ ),
    .B(\MuI._2130_ ),
    .Y(\MuI._2131_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6263_  (.A(\MuI._2131_ ),
    .B(\MuI._2104_ ),
    .Y(\MuI._2133_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6264_  (.A1(\MuI._1043_ ),
    .A2(\MuI._1285_ ),
    .A3(\MuI._2016_ ),
    .B1(\MuI._2014_ ),
    .X(\MuI._2134_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6265_  (.A_N(\MuI._2133_ ),
    .B(\MuI._2134_ ),
    .X(\MuI._2135_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6266_  (.A_N(\MuI._2134_ ),
    .B(\MuI._2133_ ),
    .X(\MuI._2136_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6267_  (.A(\MuI._2135_ ),
    .B(\MuI._2136_ ),
    .Y(\MuI._2137_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6268_  (.A(\MuI._2018_ ),
    .B(\MuI._2026_ ),
    .X(\MuI._2138_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6269_  (.A(\MuI._2137_ ),
    .B(\MuI._2138_ ),
    .X(\MuI._2139_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6270_  (.A(\MuI._2126_ ),
    .B(\MuI._2139_ ),
    .Y(\MuI._2140_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6271_  (.A(\MuI._2043_ ),
    .B_N(\MuI._2063_ ),
    .X(\MuI._2141_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6272_  (.A(\MuI._2140_ ),
    .B(\MuI._2141_ ),
    .Y(\MuI._2142_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6273_  (.A(\MuI._2108_ ),
    .B(\MuI._2142_ ),
    .Y(\MuI._2144_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6274_  (.A_N(\MuI._2107_ ),
    .B(\MuI._2144_ ),
    .X(\MuI._2145_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._6275_  (.A1(\MuI._2074_ ),
    .A2(\MuI._2101_ ),
    .B1_N(\MuI._2073_ ),
    .Y(\MuI._2146_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6276_  (.A_N(\MuI._2054_ ),
    .B(\MuI._2050_ ),
    .X(\MuI._2147_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6277_  (.A1(\MuI._2056_ ),
    .A2(\MuI._2061_ ),
    .B1(\MuI._2147_ ),
    .Y(\MuI._2148_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6278_  (.A(\MuI._2146_ ),
    .B(\MuI._2148_ ),
    .X(\MuI._2149_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6279_  (.A1(\MuI._2057_ ),
    .A2(\MuI._2060_ ),
    .B1_N(\MuI._2058_ ),
    .X(\MuI._2150_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6280_  (.A(\MuI._2149_ ),
    .B(\MuI._2150_ ),
    .X(\MuI._2151_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6281_  (.A(\MuI._2107_ ),
    .B(\MuI._2144_ ),
    .X(\MuI._2152_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6282_  (.A(\MuI._2151_ ),
    .B(\MuI._2152_ ),
    .Y(\MuI._2153_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6283_  (.A(\MuI._2145_ ),
    .B(\MuI._2153_ ),
    .Y(\MuI._2155_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6284_  (.A_N(\MuI._2140_ ),
    .B(\MuI._2141_ ),
    .X(\MuI._2156_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6285_  (.A1(\MuI._2119_ ),
    .A2(\MuI._2125_ ),
    .B1(\MuI._2117_ ),
    .Y(\MuI._2157_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6286_  (.A(\MuI._2156_ ),
    .B(\MuI._2157_ ),
    .Y(\MuI._2158_ ));
 sky130_fd_sc_hd__a32o_1 \MuI._6287_  (.A1(\MuI._2914_ ),
    .A2(\MuI._0460_ ),
    .A3(\MuI._2122_ ),
    .B1(\MuI._2120_ ),
    .B2(\MuI._2849_ ),
    .X(\MuI._2159_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6288_  (.A(\MuI._2158_ ),
    .B(\MuI._2159_ ),
    .Y(\MuI._2160_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6289_  (.A_N(\MuI._2138_ ),
    .B(\MuI._2137_ ),
    .X(\MuI._2161_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6290_  (.A(\MuI._2126_ ),
    .B(\MuI._2139_ ),
    .Y(\MuI._2162_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6291_  (.A1(\MuI._2127_ ),
    .A2(\MuI._2129_ ),
    .B1_N(\MuI._2128_ ),
    .X(\MuI._2163_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6292_  (.A(\MuI._0581_ ),
    .B(\MuI._1285_ ),
    .Y(\MuI._2164_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6293_  (.A(\MuI._2164_ ),
    .B(\MuI._1846_ ),
    .Y(\MuI._2166_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6294_  (.A(\MuI._2163_ ),
    .B(\MuI._2166_ ),
    .Y(\MuI._2167_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6295_  (.A1(\MuI._2131_ ),
    .A2(\MuI._2104_ ),
    .B1(\MuI._2135_ ),
    .Y(\MuI._2168_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6296_  (.A(\MuI._2167_ ),
    .B(\MuI._2168_ ),
    .X(\MuI._2169_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6297_  (.A(\MuI._0746_ ),
    .B(\MuI._0790_ ),
    .C(\MuI._1153_ ),
    .D(\MuI._1032_ ),
    .X(\MuI._2170_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6298_  (.A1(\MuI._0801_ ),
    .A2(\MuI._1164_ ),
    .B1(\MuI._1043_ ),
    .B2(\MuI._0746_ ),
    .Y(\MuI._2171_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6299_  (.A(\MuI._2170_ ),
    .B(\MuI._2171_ ),
    .Y(\MuI._2172_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6300_  (.A(\MuI._0878_ ),
    .B(\MuI._1494_ ),
    .C(\MuI._2172_ ),
    .X(\MuI._2173_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6301_  (.A1(\MuI._0889_ ),
    .A2(\MuI._1494_ ),
    .B1(\MuI._2172_ ),
    .Y(\MuI._2174_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6302_  (.A(\MuI._2173_ ),
    .B(\MuI._2174_ ),
    .Y(\MuI._2175_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6303_  (.A(\MuI._2109_ ),
    .B(\MuI._2113_ ),
    .Y(\MuI._2177_ ));
 sky130_fd_sc_hd__xnor2_2 \MuI._6304_  (.A(\MuI._2175_ ),
    .B(\MuI._2177_ ),
    .Y(\MuI._2178_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._6305_  (.A1(\MuI._0625_ ),
    .A2(\MuI._2077_ ),
    .B1(\MuI._3091_ ),
    .B2(\MuI._0372_ ),
    .X(\MuI._2179_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6306_  (.A1(\MuI._2077_ ),
    .A2(\MuI._2120_ ),
    .B1_N(\MuI._2179_ ),
    .X(\MuI._2180_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6307_  (.A(\MuI._2849_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._2181_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6308_  (.A(\MuI._2180_ ),
    .B(\MuI._2181_ ),
    .Y(\MuI._2182_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6309_  (.A(\MuI._2178_ ),
    .B(\MuI._2182_ ),
    .X(\MuI._2183_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6310_  (.A(\MuI._2169_ ),
    .B(\MuI._2183_ ),
    .X(\MuI._2184_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6311_  (.A1(\MuI._2161_ ),
    .A2(\MuI._2162_ ),
    .B1(\MuI._2184_ ),
    .Y(\MuI._2185_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6312_  (.A(\MuI._2161_ ),
    .B(\MuI._2162_ ),
    .C(\MuI._2184_ ),
    .X(\MuI._2186_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6313_  (.A(\MuI._2185_ ),
    .B(\MuI._2186_ ),
    .Y(\MuI._2188_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6314_  (.A(\MuI._2108_ ),
    .B_N(\MuI._2142_ ),
    .X(\MuI._2189_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6315_  (.A(\MuI._2188_ ),
    .B(\MuI._2189_ ),
    .Y(\MuI._2190_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6316_  (.A(\MuI._2160_ ),
    .B(\MuI._2190_ ),
    .Y(\MuI._2191_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6317_  (.A(\MuI._2160_ ),
    .B(\MuI._2190_ ),
    .X(\MuI._2192_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6318_  (.A(\MuI._2191_ ),
    .B(\MuI._2192_ ),
    .Y(\MuI._2193_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6319_  (.A(\MuI._2155_ ),
    .B_N(\MuI._2193_ ),
    .X(\MuI._2194_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6320_  (.A(\MuI._2193_ ),
    .B(\MuI._2155_ ),
    .X(\MuI._2195_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6321_  (.A(\MuI._2150_ ),
    .B_N(\MuI._2149_ ),
    .X(\MuI._2196_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6322_  (.A1(\MuI._2146_ ),
    .A2(\MuI._2148_ ),
    .B1(\MuI._2196_ ),
    .Y(\MuI._2197_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6323_  (.A(\MuI._2195_ ),
    .B_N(\MuI._2197_ ),
    .X(\MuI._2199_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6324_  (.A(\MuI._2157_ ),
    .B(\MuI._2140_ ),
    .C_N(\MuI._2141_ ),
    .X(\MuI._2200_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6325_  (.A(\MuI._2158_ ),
    .B(\MuI._2159_ ),
    .Y(\MuI._2201_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6326_  (.A(\MuI._2188_ ),
    .B(\MuI._2189_ ),
    .Y(\MuI._2202_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6327_  (.A(\MuI._2178_ ),
    .Y(\MuI._2203_ ));
 sky130_fd_sc_hd__o32a_1 \MuI._6328_  (.A1(\MuI._2173_ ),
    .A2(\MuI._2174_ ),
    .A3(\MuI._2177_ ),
    .B1(\MuI._2203_ ),
    .B2(\MuI._2182_ ),
    .X(\MuI._2204_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6329_  (.A(\MuI._2185_ ),
    .B(\MuI._2204_ ),
    .Y(\MuI._2205_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._6330_  (.A1_N(\MuI._2077_ ),
    .A2_N(\MuI._2120_ ),
    .B1(\MuI._2180_ ),
    .B2(\MuI._2181_ ),
    .X(\MuI._2206_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6331_  (.A(\MuI._2205_ ),
    .B(\MuI._2206_ ),
    .Y(\MuI._2207_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6332_  (.A_N(\MuI._2168_ ),
    .B(\MuI._2167_ ),
    .X(\MuI._2208_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6333_  (.A(\MuI._2169_ ),
    .B(\MuI._2183_ ),
    .Y(\MuI._2210_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6334_  (.A(\MuI._2163_ ),
    .B_N(\MuI._2166_ ),
    .X(\MuI._2211_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6335_  (.A(\MuI._1857_ ),
    .B(\MuI._1879_ ),
    .Y(\MuI._2212_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6336_  (.A(\MuI._2211_ ),
    .B(\MuI._2212_ ),
    .Y(\MuI._2213_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6337_  (.A1(\MuI._0889_ ),
    .A2(\MuI._1043_ ),
    .B1(\MuI._1945_ ),
    .Y(\MuI._2214_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6338_  (.A(\MuI._1956_ ),
    .B(\MuI._2214_ ),
    .Y(\MuI._2215_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6339_  (.A(\MuI._2170_ ),
    .B(\MuI._2173_ ),
    .Y(\MuI._2216_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6340_  (.A(\MuI._2215_ ),
    .B(\MuI._2216_ ),
    .Y(\MuI._2217_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6341_  (.A1(\MuI._0625_ ),
    .A2(\MuI._1494_ ),
    .B1(\MuI._2077_ ),
    .B2(\MuI._0372_ ),
    .Y(\MuI._2218_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6342_  (.A(\MuI._0372_ ),
    .B(\MuI._0625_ ),
    .C(\MuI._1494_ ),
    .D(\MuI._2077_ ),
    .X(\MuI._2219_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6343_  (.A(\MuI._2218_ ),
    .B(\MuI._2219_ ),
    .X(\MuI._2221_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6344_  (.A(\MuI._3091_ ),
    .B(\MuI._0460_ ),
    .Y(\MuI._2222_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6345_  (.A(\MuI._2221_ ),
    .B(\MuI._2222_ ),
    .X(\MuI._2223_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6346_  (.A(\MuI._2217_ ),
    .B(\MuI._2223_ ),
    .Y(\MuI._2224_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6347_  (.A(\MuI._2217_ ),
    .B(\MuI._2223_ ),
    .X(\MuI._2225_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6348_  (.A(\MuI._2224_ ),
    .B(\MuI._2225_ ),
    .Y(\MuI._2226_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6349_  (.A(\MuI._2213_ ),
    .B(\MuI._2226_ ),
    .Y(\MuI._2227_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6350_  (.A1(\MuI._2208_ ),
    .A2(\MuI._2210_ ),
    .B1_N(\MuI._2227_ ),
    .X(\MuI._2228_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6351_  (.A(\MuI._2208_ ),
    .B(\MuI._2210_ ),
    .C_N(\MuI._2227_ ),
    .X(\MuI._2229_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6352_  (.A(\MuI._2228_ ),
    .B_N(\MuI._2229_ ),
    .X(\MuI._2230_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6353_  (.A(\MuI._2207_ ),
    .B(\MuI._2230_ ),
    .Y(\MuI._2232_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6354_  (.A(\MuI._2207_ ),
    .B(\MuI._2230_ ),
    .X(\MuI._2233_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6355_  (.A(\MuI._2232_ ),
    .B(\MuI._2233_ ),
    .Y(\MuI._2234_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6356_  (.A1(\MuI._2202_ ),
    .A2(\MuI._2191_ ),
    .B1(\MuI._2234_ ),
    .X(\MuI._2235_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6357_  (.A(\MuI._2234_ ),
    .B(\MuI._2202_ ),
    .C(\MuI._2191_ ),
    .Y(\MuI._2236_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._6358_  (.A1(\MuI._2200_ ),
    .A2(\MuI._2201_ ),
    .B1(\MuI._2235_ ),
    .C1(\MuI._2236_ ),
    .Y(\MuI._2237_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6359_  (.A1(\MuI._2235_ ),
    .A2(\MuI._2236_ ),
    .B1(\MuI._2200_ ),
    .C1(\MuI._2201_ ),
    .X(\MuI._2238_ ));
 sky130_fd_sc_hd__a211oi_1 \MuI._6360_  (.A1(\MuI._2194_ ),
    .A2(\MuI._2199_ ),
    .B1(\MuI._2237_ ),
    .C1(\MuI._2238_ ),
    .Y(\MuI._2239_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6361_  (.A1(\MuI._2237_ ),
    .A2(\MuI._2238_ ),
    .B1(\MuI._2194_ ),
    .C1(\MuI._2199_ ),
    .X(\MuI._2240_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6362_  (.A(\MuI._2239_ ),
    .B(\MuI._2240_ ),
    .X(\MuI._2241_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6363_  (.A(\MuI._2197_ ),
    .B(\MuI._2195_ ),
    .X(\MuI._2243_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6364_  (.A1(\MuI._2102_ ),
    .A2(\MuI._2103_ ),
    .B1(\MuI._2106_ ),
    .X(\MuI._2244_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6365_  (.A(\MuI._1930_ ),
    .B_N(\MuI._1936_ ),
    .X(\MuI._2245_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6366_  (.A(\MuI._1929_ ),
    .B(\MuI._1937_ ),
    .Y(\MuI._2246_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6367_  (.A(\MuI._2081_ ),
    .B(\MuI._2076_ ),
    .C(\MuI._2080_ ),
    .X(\MuI._2247_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6368_  (.A1(\MuI._2081_ ),
    .A2(\MuI._2080_ ),
    .B1(\MuI._2076_ ),
    .Y(\MuI._2248_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6369_  (.A(\MuI._2247_ ),
    .B(\MuI._2248_ ),
    .X(\MuI._2249_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6370_  (.A1(\MuI._2245_ ),
    .A2(\MuI._2246_ ),
    .B1(\MuI._2249_ ),
    .Y(\MuI._2250_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6371_  (.A(\MuI._2250_ ),
    .Y(\MuI._2251_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6372_  (.A(\MuI._2245_ ),
    .B(\MuI._2246_ ),
    .C(\MuI._2249_ ),
    .X(\MuI._2252_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._6373_  (.A1_N(\MuI._0867_ ),
    .A2_N(\MuI._2682_ ),
    .B1(\MuI._2087_ ),
    .B2(\MuI._2089_ ),
    .X(\MuI._2254_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6374_  (.A(\MuI._2090_ ),
    .B(\MuI._2254_ ),
    .Y(\MuI._2255_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6375_  (.A1(\MuI._1942_ ),
    .A2(\MuI._1944_ ),
    .B1_N(\MuI._1943_ ),
    .X(\MuI._2256_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6376_  (.A(\MuI._2255_ ),
    .B(\MuI._2256_ ),
    .Y(\MuI._2257_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6377_  (.A1(\MuI._0603_ ),
    .A2(\MuI._2594_ ),
    .B1(\MuI._2797_ ),
    .B2(\MuI._2826_ ),
    .Y(\MuI._2258_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6378_  (.A(\MuI._2826_ ),
    .B(\MuI._0603_ ),
    .C(\MuI._2594_ ),
    .D(\MuI._2797_ ),
    .X(\MuI._2259_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6379_  (.A(\MuI._2258_ ),
    .B(\MuI._2259_ ),
    .Y(\MuI._2260_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6380_  (.A(\MuI._2789_ ),
    .B(\MuI._0438_ ),
    .Y(\MuI._2261_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6381_  (.A(\MuI._2260_ ),
    .B(\MuI._2261_ ),
    .Y(\MuI._2262_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6382_  (.A(\MuI._2257_ ),
    .B(\MuI._2262_ ),
    .Y(\MuI._2263_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6383_  (.A(\MuI._2257_ ),
    .B(\MuI._2262_ ),
    .X(\MuI._2265_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6384_  (.A(\MuI._2263_ ),
    .B(\MuI._2265_ ),
    .Y(\MuI._2266_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6385_  (.A(\MuI._2250_ ),
    .B(\MuI._2252_ ),
    .C(\MuI._2266_ ),
    .X(\MuI._2267_ ));
 sky130_fd_sc_hd__nand3b_1 \MuI._6386_  (.A_N(\MuI._1887_ ),
    .B(\MuI._2851_ ),
    .C(\MuI._0526_ ),
    .Y(\MuI._2268_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6387_  (.A(\MuI._2065_ ),
    .B(\MuI._2268_ ),
    .X(\MuI._2269_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6388_  (.A1(\MuI._2083_ ),
    .A2(\MuI._2084_ ),
    .B1(\MuI._2098_ ),
    .Y(\MuI._2270_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6389_  (.A(\MuI._1966_ ),
    .B(\MuI._1969_ ),
    .X(\MuI._2271_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6390_  (.A(\MuI._1966_ ),
    .B(\MuI._1969_ ),
    .X(\MuI._2272_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6391_  (.A1(\MuI._2271_ ),
    .A2(\MuI._1975_ ),
    .B1(\MuI._2272_ ),
    .X(\MuI._2273_ ));
 sky130_fd_sc_hd__and4b_1 \MuI._6392_  (.A_N(\MuI._2269_ ),
    .B(\MuI._2270_ ),
    .C(\MuI._2100_ ),
    .D(\MuI._2273_ ),
    .X(\MuI._2274_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6393_  (.A1(\MuI._2271_ ),
    .A2(\MuI._1975_ ),
    .B1(\MuI._2272_ ),
    .Y(\MuI._2276_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._6394_  (.A1_N(\MuI._2100_ ),
    .A2_N(\MuI._2270_ ),
    .B1(\MuI._2269_ ),
    .B2(\MuI._2276_ ),
    .X(\MuI._2277_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6395_  (.A1(\MuI._2251_ ),
    .A2(\MuI._2267_ ),
    .B1(\MuI._2274_ ),
    .C1(\MuI._2277_ ),
    .X(\MuI._2278_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._6396_  (.A1(\MuI._2274_ ),
    .A2(\MuI._2277_ ),
    .B1(\MuI._2251_ ),
    .C1(\MuI._2267_ ),
    .Y(\MuI._2279_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6397_  (.A(\MuI._2067_ ),
    .B(\MuI._2070_ ),
    .Y(\MuI._2280_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6398_  (.A(\MuI._2071_ ),
    .B(\MuI._2280_ ),
    .Y(\MuI._2281_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6399_  (.A(\MuI._2278_ ),
    .B(\MuI._2279_ ),
    .C(\MuI._2281_ ),
    .X(\MuI._2282_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6400_  (.A(\MuI._2107_ ),
    .B(\MuI._2244_ ),
    .C(\MuI._2282_ ),
    .X(\MuI._2283_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6401_  (.A(\MuI._2100_ ),
    .B(\MuI._2270_ ),
    .Y(\MuI._2284_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6402_  (.A(\MuI._2276_ ),
    .B(\MuI._2269_ ),
    .C(\MuI._2284_ ),
    .X(\MuI._2285_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6403_  (.A(\MuI._2092_ ),
    .B(\MuI._2097_ ),
    .Y(\MuI._2287_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6404_  (.A1(\MuI._2053_ ),
    .A2(\MuI._2085_ ),
    .A3(\MuI._2091_ ),
    .B1(\MuI._2287_ ),
    .X(\MuI._2288_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6405_  (.A1(\MuI._2285_ ),
    .A2(\MuI._2278_ ),
    .B1(\MuI._2288_ ),
    .X(\MuI._2289_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6406_  (.A(\MuI._2285_ ),
    .B(\MuI._2278_ ),
    .C(\MuI._2288_ ),
    .Y(\MuI._2290_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6407_  (.A(\MuI._2289_ ),
    .B(\MuI._2290_ ),
    .X(\MuI._2291_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6408_  (.A1(\MuI._2093_ ),
    .A2(\MuI._2096_ ),
    .B1_N(\MuI._2094_ ),
    .X(\MuI._2292_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6409_  (.A(\MuI._2291_ ),
    .B(\MuI._2292_ ),
    .X(\MuI._2293_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6410_  (.A1(\MuI._2107_ ),
    .A2(\MuI._2244_ ),
    .B1(\MuI._2282_ ),
    .Y(\MuI._2294_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6411_  (.A(\MuI._2283_ ),
    .B(\MuI._2293_ ),
    .C(\MuI._2294_ ),
    .Y(\MuI._2295_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6412_  (.A(\MuI._2283_ ),
    .B(\MuI._2295_ ),
    .Y(\MuI._2296_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6413_  (.A(\MuI._2151_ ),
    .B(\MuI._2152_ ),
    .X(\MuI._2298_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6414_  (.A(\MuI._2153_ ),
    .B(\MuI._2298_ ),
    .Y(\MuI._2299_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6415_  (.A_N(\MuI._2296_ ),
    .B(\MuI._2299_ ),
    .X(\MuI._2300_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6416_  (.A(\MuI._2299_ ),
    .B(\MuI._2296_ ),
    .X(\MuI._2301_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6417_  (.A(\MuI._2292_ ),
    .B_N(\MuI._2291_ ),
    .X(\MuI._2302_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6418_  (.A(\MuI._2289_ ),
    .B(\MuI._2302_ ),
    .Y(\MuI._2303_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6419_  (.A_N(\MuI._2301_ ),
    .B(\MuI._2303_ ),
    .X(\MuI._2304_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6420_  (.A(\MuI._2300_ ),
    .B(\MuI._2304_ ),
    .Y(\MuI._2305_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6421_  (.A(\MuI._2243_ ),
    .B(\MuI._2305_ ),
    .Y(\MuI._2306_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6422_  (.A(\MuI._2241_ ),
    .B(\MuI._2306_ ),
    .X(\MuI._2307_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6423_  (.A(\MuI._2303_ ),
    .B(\MuI._2301_ ),
    .Y(\MuI._2309_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6424_  (.A1(\MuI._2278_ ),
    .A2(\MuI._2279_ ),
    .B1(\MuI._2281_ ),
    .Y(\MuI._2310_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6425_  (.A(\MuI._1941_ ),
    .B(\MuI._1955_ ),
    .X(\MuI._2311_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6426_  (.A1(\MuI._2250_ ),
    .A2(\MuI._2252_ ),
    .B1(\MuI._2266_ ),
    .Y(\MuI._2312_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6427_  (.A(\MuI._1977_ ),
    .B(\MuI._2267_ ),
    .C(\MuI._2312_ ),
    .X(\MuI._2313_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6428_  (.A1(\MuI._2267_ ),
    .A2(\MuI._2312_ ),
    .B1(\MuI._1977_ ),
    .Y(\MuI._2314_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._6429_  (.A1(\MuI._1939_ ),
    .A2(\MuI._2311_ ),
    .B1(\MuI._2313_ ),
    .C1(\MuI._2314_ ),
    .Y(\MuI._2315_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6430_  (.A1(\MuI._2313_ ),
    .A2(\MuI._2314_ ),
    .B1(\MuI._1939_ ),
    .C1(\MuI._2311_ ),
    .X(\MuI._2316_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6431_  (.A(\MuI._2276_ ),
    .B(\MuI._2269_ ),
    .Y(\MuI._2317_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6432_  (.A(\MuI._2315_ ),
    .B(\MuI._2316_ ),
    .C(\MuI._2317_ ),
    .X(\MuI._2318_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6433_  (.A(\MuI._2282_ ),
    .B(\MuI._2310_ ),
    .C(\MuI._2318_ ),
    .X(\MuI._2320_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6434_  (.A1(\MuI._2090_ ),
    .A2(\MuI._2254_ ),
    .A3(\MuI._2256_ ),
    .B1(\MuI._2263_ ),
    .X(\MuI._2321_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6435_  (.A1(\MuI._2313_ ),
    .A2(\MuI._2315_ ),
    .B1_N(\MuI._2321_ ),
    .X(\MuI._2322_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6436_  (.A(\MuI._2313_ ),
    .B(\MuI._2315_ ),
    .C_N(\MuI._2321_ ),
    .X(\MuI._2323_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6437_  (.A_N(\MuI._2322_ ),
    .B(\MuI._2323_ ),
    .X(\MuI._2324_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6438_  (.A1(\MuI._2258_ ),
    .A2(\MuI._2261_ ),
    .B1_N(\MuI._2259_ ),
    .X(\MuI._2325_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6439_  (.A(\MuI._2324_ ),
    .B(\MuI._2325_ ),
    .Y(\MuI._2326_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6440_  (.A1(\MuI._2282_ ),
    .A2(\MuI._2310_ ),
    .B1(\MuI._2318_ ),
    .Y(\MuI._2327_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6441_  (.A(\MuI._2320_ ),
    .B(\MuI._2326_ ),
    .C(\MuI._2327_ ),
    .Y(\MuI._2328_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6442_  (.A1(\MuI._2283_ ),
    .A2(\MuI._2294_ ),
    .B1(\MuI._2293_ ),
    .X(\MuI._2329_ ));
 sky130_fd_sc_hd__a211oi_2 \MuI._6443_  (.A1(\MuI._2320_ ),
    .A2(\MuI._2328_ ),
    .B1(\MuI._2295_ ),
    .C1(\MuI._2329_ ),
    .Y(\MuI._2331_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6444_  (.A(\MuI._2325_ ),
    .Y(\MuI._2332_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6445_  (.A1(\MuI._2324_ ),
    .A2(\MuI._2332_ ),
    .B1(\MuI._2322_ ),
    .X(\MuI._2333_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._6446_  (.A1(\MuI._2295_ ),
    .A2(\MuI._2329_ ),
    .B1(\MuI._2320_ ),
    .C1(\MuI._2328_ ),
    .Y(\MuI._2334_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6447_  (.A_N(\MuI._2331_ ),
    .B(\MuI._2334_ ),
    .X(\MuI._2335_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6448_  (.A(\MuI._2333_ ),
    .B(\MuI._2335_ ),
    .X(\MuI._2336_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6449_  (.A(\MuI._2309_ ),
    .B(\MuI._2331_ ),
    .C(\MuI._2336_ ),
    .Y(\MuI._2337_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6450_  (.A1(\MuI._2331_ ),
    .A2(\MuI._2336_ ),
    .B1(\MuI._2309_ ),
    .X(\MuI._2338_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6451_  (.A(\MuI._2337_ ),
    .B(\MuI._2338_ ),
    .X(\MuI._2339_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6452_  (.A(\MuI._2333_ ),
    .B(\MuI._2335_ ),
    .Y(\MuI._2340_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6453_  (.A_N(\MuI._1957_ ),
    .B(\MuI._1926_ ),
    .X(\MuI._2342_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6454_  (.A1(\MuI._1958_ ),
    .A2(\MuI._1961_ ),
    .B1(\MuI._2342_ ),
    .Y(\MuI._2343_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6455_  (.A_N(\MuI._1948_ ),
    .B(\MuI._1947_ ),
    .X(\MuI._2344_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6456_  (.A1(\MuI._1949_ ),
    .A2(\MuI._1954_ ),
    .B1(\MuI._2344_ ),
    .Y(\MuI._2345_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6457_  (.A1(\MuI._1950_ ),
    .A2(\MuI._1953_ ),
    .B1_N(\MuI._1951_ ),
    .X(\MuI._2346_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6458_  (.A(\MuI._2343_ ),
    .B(\MuI._2345_ ),
    .X(\MuI._2347_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6459_  (.A(\MuI._2346_ ),
    .B_N(\MuI._2347_ ),
    .X(\MuI._2348_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6460_  (.A1(\MuI._2343_ ),
    .A2(\MuI._2345_ ),
    .B1(\MuI._2348_ ),
    .Y(\MuI._2349_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6461_  (.A(\MuI._2320_ ),
    .B(\MuI._2327_ ),
    .Y(\MuI._2350_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6462_  (.A(\MuI._2326_ ),
    .B(\MuI._2350_ ),
    .Y(\MuI._2351_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6463_  (.A(\MuI._2347_ ),
    .B(\MuI._2346_ ),
    .X(\MuI._2353_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6464_  (.A(\MuI._1962_ ),
    .B_N(\MuI._1980_ ),
    .X(\MuI._2354_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6465_  (.A1(\MuI._2315_ ),
    .A2(\MuI._2316_ ),
    .B1(\MuI._2317_ ),
    .Y(\MuI._2355_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6466_  (.A(\MuI._2318_ ),
    .B(\MuI._2355_ ),
    .Y(\MuI._2356_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6467_  (.A(\MuI._2354_ ),
    .B(\MuI._2356_ ),
    .Y(\MuI._2357_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6468_  (.A(\MuI._2354_ ),
    .B(\MuI._2356_ ),
    .Y(\MuI._2358_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6469_  (.A1(\MuI._2353_ ),
    .A2(\MuI._2357_ ),
    .B1_N(\MuI._2358_ ),
    .X(\MuI._2359_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6470_  (.A(\MuI._2351_ ),
    .B(\MuI._2359_ ),
    .Y(\MuI._2360_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6471_  (.A_N(\MuI._2359_ ),
    .B(\MuI._2351_ ),
    .X(\MuI._2361_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6472_  (.A1(\MuI._2349_ ),
    .A2(\MuI._2360_ ),
    .B1(\MuI._2361_ ),
    .Y(\MuI._2362_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6473_  (.A(\MuI._2340_ ),
    .B(\MuI._2362_ ),
    .Y(\MuI._2364_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6474_  (.A(\MuI._2340_ ),
    .B(\MuI._2362_ ),
    .X(\MuI._2365_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6475_  (.A(\MuI._2364_ ),
    .B(\MuI._2365_ ),
    .X(\MuI._2366_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6476_  (.A(\MuI._2307_ ),
    .B(\MuI._2339_ ),
    .C(\MuI._2366_ ),
    .X(\MuI._2367_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6477_  (.A(\MuI._2353_ ),
    .B(\MuI._2357_ ),
    .Y(\MuI._2368_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6478_  (.A_N(\MuI._1983_ ),
    .B(\MuI._1981_ ),
    .X(\MuI._2369_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6479_  (.A1(\MuI._1924_ ),
    .A2(\MuI._1984_ ),
    .B1(\MuI._2369_ ),
    .Y(\MuI._2370_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6480_  (.A(\MuI._2368_ ),
    .B(\MuI._2370_ ),
    .X(\MuI._2371_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6481_  (.A(\MuI._2368_ ),
    .B(\MuI._2370_ ),
    .Y(\MuI._2372_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6482_  (.A(\MuI._1922_ ),
    .B_N(\MuI._1921_ ),
    .X(\MuI._2373_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._6483_  (.A1(\MuI._1919_ ),
    .A2(\MuI._1920_ ),
    .B1(\MuI._2373_ ),
    .Y(\MuI._2375_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6484_  (.A(\MuI._2372_ ),
    .B_N(\MuI._2375_ ),
    .X(\MuI._2376_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6485_  (.A(\MuI._2349_ ),
    .B(\MuI._2360_ ),
    .Y(\MuI._2377_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6486_  (.A1(\MuI._2371_ ),
    .A2(\MuI._2376_ ),
    .B1(\MuI._2377_ ),
    .Y(\MuI._2378_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6487_  (.A(\MuI._2377_ ),
    .B(\MuI._2371_ ),
    .C(\MuI._2376_ ),
    .X(\MuI._2379_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6488_  (.A(\MuI._2378_ ),
    .B(\MuI._2379_ ),
    .Y(\MuI._2380_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6489_  (.A(\MuI._2375_ ),
    .B(\MuI._2372_ ),
    .X(\MuI._2381_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6490_  (.A1(\MuI._1917_ ),
    .A2(\MuI._1992_ ),
    .B1(\MuI._1990_ ),
    .Y(\MuI._2382_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6491_  (.A(\MuI._2381_ ),
    .B(\MuI._2382_ ),
    .X(\MuI._2383_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6492_  (.A(\MuI._2380_ ),
    .B(\MuI._2383_ ),
    .Y(\MuI._2384_ ));
 sky130_fd_sc_hd__a2111o_1 \MuI._6493_  (.A1(\MuI._0793_ ),
    .A2(\MuI._1841_ ),
    .B1(\MuI._2005_ ),
    .C1(\MuI._2367_ ),
    .D1(\MuI._2384_ ),
    .X(\MuI._2386_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6494_  (.A(\MuI._2338_ ),
    .B(\MuI._2364_ ),
    .Y(\MuI._2387_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6495_  (.A(\MuI._2307_ ),
    .B(\MuI._2337_ ),
    .C(\MuI._2387_ ),
    .X(\MuI._2388_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6496_  (.A(\MuI._2243_ ),
    .B(\MuI._2305_ ),
    .X(\MuI._2389_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6497_  (.A1(\MuI._2240_ ),
    .A2(\MuI._2389_ ),
    .B1_N(\MuI._2239_ ),
    .X(\MuI._2390_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6498_  (.A(\MuI._2381_ ),
    .B(\MuI._2382_ ),
    .Y(\MuI._2391_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6499_  (.A1(\MuI._2378_ ),
    .A2(\MuI._2391_ ),
    .B1_N(\MuI._2379_ ),
    .Y(\MuI._2392_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6500_  (.A1(\MuI._1909_ ),
    .A2(\MuI._1915_ ),
    .B1(\MuI._1993_ ),
    .X(\MuI._2393_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6501_  (.A1(\MuI._2393_ ),
    .A2(\MuI._2001_ ),
    .B1(\MuI._1995_ ),
    .Y(\MuI._2394_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6502_  (.A(\MuI._2384_ ),
    .B_N(\MuI._2394_ ),
    .X(\MuI._2395_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6503_  (.A1(\MuI._2392_ ),
    .A2(\MuI._2395_ ),
    .B1(\MuI._2367_ ),
    .X(\MuI._2397_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6504_  (.A(\MuI._2388_ ),
    .B(\MuI._2390_ ),
    .C(\MuI._2397_ ),
    .X(\MuI._2398_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6505_  (.A(\MuI._2231_ ),
    .B(\MuI._2253_ ),
    .Y(\MuI._2399_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6506_  (.A1(\MuI._2044_ ),
    .A2(\MuI._2088_ ),
    .B1_N(\MuI._2033_ ),
    .X(\MuI._2400_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6507_  (.A(\MuI._2211_ ),
    .B(\MuI._2212_ ),
    .Y(\MuI._2401_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6508_  (.A(\MuI._2213_ ),
    .B(\MuI._2226_ ),
    .Y(\MuI._2402_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6509_  (.A(\MuI._1912_ ),
    .B(\MuI._2110_ ),
    .X(\MuI._2403_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6510_  (.A(\MuI._2121_ ),
    .B(\MuI._2403_ ),
    .Y(\MuI._2404_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6511_  (.A1(\MuI._2401_ ),
    .A2(\MuI._2402_ ),
    .B1(\MuI._2404_ ),
    .X(\MuI._2405_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6512_  (.A1(\MuI._2000_ ),
    .A2(\MuI._2099_ ),
    .B1(\MuI._1989_ ),
    .Y(\MuI._2406_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6513_  (.A(\MuI._2405_ ),
    .B(\MuI._2406_ ),
    .Y(\MuI._2408_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6514_  (.A_N(\MuI._2400_ ),
    .B(\MuI._2408_ ),
    .X(\MuI._2409_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6515_  (.A_N(\MuI._2408_ ),
    .B(\MuI._2400_ ),
    .X(\MuI._2410_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6516_  (.A(\MuI._2409_ ),
    .B(\MuI._2410_ ),
    .X(\MuI._2411_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6517_  (.A_N(\MuI._2132_ ),
    .B(\MuI._1780_ ),
    .X(\MuI._2412_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6518_  (.A(\MuI._2143_ ),
    .B(\MuI._2412_ ),
    .X(\MuI._2413_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6519_  (.A(\MuI._2411_ ),
    .B(\MuI._2413_ ),
    .Y(\MuI._2414_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6520_  (.A(\MuI._2264_ ),
    .B(\MuI._2399_ ),
    .C_N(\MuI._2414_ ),
    .X(\MuI._2415_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6521_  (.A_N(\MuI._2406_ ),
    .B(\MuI._2405_ ),
    .X(\MuI._2416_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6522_  (.A1(\MuI._2264_ ),
    .A2(\MuI._2399_ ),
    .B1_N(\MuI._2414_ ),
    .Y(\MuI._2417_ ));
 sky130_fd_sc_hd__o211ai_1 \MuI._6523_  (.A1(\MuI._2416_ ),
    .A2(\MuI._2409_ ),
    .B1(\MuI._2415_ ),
    .C1(\MuI._2417_ ),
    .Y(\MuI._2419_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6524_  (.A(\MuI._2209_ ),
    .B(\MuI._2275_ ),
    .Y(\MuI._2420_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6525_  (.A1(\MuI._2415_ ),
    .A2(\MuI._2419_ ),
    .B1(\MuI._2420_ ),
    .X(\MuI._2421_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6526_  (.A(\MuI._2420_ ),
    .B(\MuI._2415_ ),
    .C(\MuI._2419_ ),
    .X(\MuI._2422_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6527_  (.A(\MuI._2422_ ),
    .Y(\MuI._2423_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6528_  (.A(\MuI._2421_ ),
    .B(\MuI._2423_ ),
    .Y(\MuI._2424_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6529_  (.A1(\MuI._2415_ ),
    .A2(\MuI._2417_ ),
    .B1(\MuI._2416_ ),
    .C1(\MuI._2409_ ),
    .X(\MuI._2425_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6530_  (.A(\MuI._2419_ ),
    .B(\MuI._2425_ ),
    .X(\MuI._2426_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6531_  (.A(\MuI._2411_ ),
    .B(\MuI._2413_ ),
    .X(\MuI._2427_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6532_  (.A1(\MuI._1956_ ),
    .A2(\MuI._2214_ ),
    .A3(\MuI._2216_ ),
    .B1(\MuI._2224_ ),
    .X(\MuI._2428_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6533_  (.A(\MuI._2228_ ),
    .B(\MuI._2428_ ),
    .Y(\MuI._2430_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6534_  (.A1(\MuI._2221_ ),
    .A2(\MuI._2222_ ),
    .B1_N(\MuI._2219_ ),
    .Y(\MuI._2431_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6535_  (.A(\MuI._2430_ ),
    .B(\MuI._2431_ ),
    .X(\MuI._2432_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6536_  (.A(\MuI._2430_ ),
    .B(\MuI._2431_ ),
    .Y(\MuI._2433_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6537_  (.A(\MuI._2432_ ),
    .B(\MuI._2433_ ),
    .Y(\MuI._2434_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6538_  (.A(\MuI._2401_ ),
    .B(\MuI._2402_ ),
    .C(\MuI._2404_ ),
    .Y(\MuI._2435_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6539_  (.A(\MuI._2405_ ),
    .B(\MuI._2435_ ),
    .Y(\MuI._2436_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6540_  (.A(\MuI._2434_ ),
    .B(\MuI._2436_ ),
    .X(\MuI._2437_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6541_  (.A(\MuI._2414_ ),
    .B(\MuI._2427_ ),
    .C_N(\MuI._2437_ ),
    .X(\MuI._2438_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6542_  (.A_N(\MuI._2428_ ),
    .B(\MuI._2228_ ),
    .X(\MuI._2439_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6543_  (.A1(\MuI._2414_ ),
    .A2(\MuI._2427_ ),
    .B1_N(\MuI._2437_ ),
    .Y(\MuI._2441_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._6544_  (.A1(\MuI._2439_ ),
    .A2(\MuI._2432_ ),
    .B1(\MuI._2438_ ),
    .C1(\MuI._2441_ ),
    .Y(\MuI._2442_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6545_  (.A(\MuI._2438_ ),
    .B(\MuI._2442_ ),
    .Y(\MuI._2443_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6546_  (.A(\MuI._2426_ ),
    .B(\MuI._2443_ ),
    .Y(\MuI._2444_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6547_  (.A(\MuI._2424_ ),
    .B(\MuI._2444_ ),
    .Y(\MuI._2445_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6548_  (.A1(\MuI._2438_ ),
    .A2(\MuI._2441_ ),
    .B1(\MuI._2439_ ),
    .C1(\MuI._2432_ ),
    .X(\MuI._2446_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6549_  (.A(\MuI._2434_ ),
    .B(\MuI._2436_ ),
    .Y(\MuI._2447_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6550_  (.A(\MuI._2437_ ),
    .B(\MuI._2447_ ),
    .Y(\MuI._2448_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6551_  (.A(\MuI._2232_ ),
    .B(\MuI._2448_ ),
    .X(\MuI._2449_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6552_  (.A(\MuI._2185_ ),
    .B(\MuI._2204_ ),
    .X(\MuI._2450_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6553_  (.A1(\MuI._2205_ ),
    .A2(\MuI._2206_ ),
    .B1(\MuI._2450_ ),
    .Y(\MuI._2452_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6554_  (.A(\MuI._2232_ ),
    .B(\MuI._2448_ ),
    .Y(\MuI._2453_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6555_  (.A(\MuI._2449_ ),
    .B(\MuI._2453_ ),
    .Y(\MuI._2454_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6556_  (.A(\MuI._2452_ ),
    .B(\MuI._2454_ ),
    .X(\MuI._2455_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6557_  (.A1(\MuI._2442_ ),
    .A2(\MuI._2446_ ),
    .B1(\MuI._2449_ ),
    .C1(\MuI._2455_ ),
    .X(\MuI._2456_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6558_  (.A(\MuI._2456_ ),
    .Y(\MuI._2457_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6559_  (.A1(\MuI._2449_ ),
    .A2(\MuI._2455_ ),
    .B1(\MuI._2442_ ),
    .C1(\MuI._2446_ ),
    .X(\MuI._2458_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6560_  (.A(\MuI._2457_ ),
    .B(\MuI._2458_ ),
    .Y(\MuI._2459_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6561_  (.A(\MuI._2445_ ),
    .B(\MuI._2459_ ),
    .Y(\MuI._2460_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6562_  (.A(\MuI._2452_ ),
    .B(\MuI._2454_ ),
    .Y(\MuI._2461_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6563_  (.A(\MuI._2235_ ),
    .B(\MuI._2237_ ),
    .Y(\MuI._2463_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6564_  (.A(\MuI._2461_ ),
    .B(\MuI._2463_ ),
    .Y(\MuI._2464_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6565_  (.A(\MuI._2461_ ),
    .B(\MuI._2463_ ),
    .X(\MuI._2465_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6566_  (.A(\MuI._2464_ ),
    .B(\MuI._2465_ ),
    .X(\MuI._2466_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6567_  (.A1(\MuI._2386_ ),
    .A2(\MuI._2398_ ),
    .B1(\MuI._2460_ ),
    .C1(\MuI._2466_ ),
    .X(\MuI._2467_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6568_  (.A(\MuI._2426_ ),
    .B(\MuI._2443_ ),
    .Y(\MuI._2468_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6569_  (.A1(\MuI._2464_ ),
    .A2(\MuI._2458_ ),
    .B1(\MuI._2456_ ),
    .X(\MuI._2469_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6570_  (.A(\MuI._2445_ ),
    .B(\MuI._2469_ ),
    .Y(\MuI._2470_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6571_  (.A1(\MuI._2422_ ),
    .A2(\MuI._2468_ ),
    .B1(\MuI._2470_ ),
    .C1(\MuI._2421_ ),
    .X(\MuI._2471_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6572_  (.A(\MuI._1758_ ),
    .B(\MuI._2297_ ),
    .X(\MuI._2472_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6573_  (.A(\MuI._2308_ ),
    .B(\MuI._2472_ ),
    .X(\MuI._2474_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6574_  (.A1(\MuI._2467_ ),
    .A2(\MuI._2471_ ),
    .B1(\MuI._2474_ ),
    .Y(\MuI._2475_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6575_  (.A(\MuI._1648_ ),
    .B(\MuI._1714_ ),
    .C(\MuI._1736_ ),
    .X(\MuI._2476_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6576_  (.A(\MuI._2476_ ),
    .Y(\MuI._2477_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6577_  (.A(\MuI._0680_ ),
    .B(\MuI._0713_ ),
    .Y(\MuI._2478_ ));
 sky130_fd_sc_hd__and4b_1 \MuI._6578_  (.A_N(\MuI._0548_ ),
    .B(\MuI._2478_ ),
    .C(\MuI._0988_ ),
    .D(\MuI._0691_ ),
    .X(\MuI._2479_ ));
 sky130_fd_sc_hd__o2bb2a_1 \MuI._6579_  (.A1_N(\MuI._2478_ ),
    .A2_N(\MuI._0988_ ),
    .B1(\MuI._0394_ ),
    .B2(\MuI._0548_ ),
    .X(\MuI._2480_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6580_  (.A(\MuI._2479_ ),
    .B(\MuI._2480_ ),
    .X(\MuI._2481_ ));
 sky130_fd_sc_hd__o311a_2 \MuI._6581_  (.A1(\MuI._1747_ ),
    .A2(\MuI._2308_ ),
    .A3(\MuI._2475_ ),
    .B1(\MuI._2477_ ),
    .C1(\MuI._2481_ ),
    .X(\MuI._2482_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6582_  (.A1(\MuI._0691_ ),
    .A2(\MuI._2478_ ),
    .B1(\MuI._0548_ ),
    .Y(\MuI._2483_ ));
 sky130_fd_sc_hd__or3_2 \MuI._6583_  (.A(\MuI._0999_ ),
    .B(\MuI._2482_ ),
    .C(\MuI._2483_ ),
    .X(\MuI._2485_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._6584_  (.A(\MuI._2485_ ),
    .X(\MuI._2486_ ));
 sky130_fd_sc_hd__clkbuf_4 \MuI._6585_  (.A(\MuI._2486_ ),
    .X(\MuI._2487_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6586_  (.A1(\MuI._0295_ ),
    .A2(\MuI._0317_ ),
    .B1(\MuI._2487_ ),
    .C1(\MuI.a_operand[23] ),
    .X(\MuI._2488_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6587_  (.A(\MuI.a_operand[23] ),
    .B(\MuI._2486_ ),
    .Y(\MuI._2489_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6588_  (.A1(\MuI.a_operand[23] ),
    .A2(\MuI._2487_ ),
    .B1(\MuI._0317_ ),
    .C1(\MuI._0295_ ),
    .X(\MuI._2490_ ));
 sky130_fd_sc_hd__a31o_1 \MuI._6589_  (.A1(\MuI.b_operand[23] ),
    .A2(\MuI._2488_ ),
    .A3(\MuI._2489_ ),
    .B1(\MuI._2490_ ),
    .X(\MuI._2491_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6590_  (.A_N(\MuI._0295_ ),
    .B(\MuI._0284_ ),
    .C(\MuI._0262_ ),
    .X(\MuI._2492_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6591_  (.A1(\MuI._0306_ ),
    .A2(\MuI._2491_ ),
    .B1(\MuI._2492_ ),
    .X(\MuI._2493_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6592_  (.A_N(\MuI._0262_ ),
    .B(\MuI._0251_ ),
    .C(\MuI._0229_ ),
    .X(\MuI._2494_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6593_  (.A1(\MuI._0273_ ),
    .A2(\MuI._2493_ ),
    .B1(\MuI._2494_ ),
    .X(\MuI._2496_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6594_  (.A_N(\MuI._0229_ ),
    .B(\MuI._0218_ ),
    .C(\MuI._0196_ ),
    .X(\MuI._2497_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6595_  (.A1(\MuI._0240_ ),
    .A2(\MuI._2496_ ),
    .B1(\MuI._2497_ ),
    .X(\MuI._2498_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6596_  (.A_N(\MuI._0196_ ),
    .B(\MuI._0185_ ),
    .C(\MuI._0163_ ),
    .X(\MuI._2499_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6597_  (.A1(\MuI._0207_ ),
    .A2(\MuI._2498_ ),
    .B1(\MuI._2499_ ),
    .X(\MuI._2500_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6598_  (.A_N(\MuI._0163_ ),
    .B(\MuI._0152_ ),
    .C(\MuI._0108_ ),
    .X(\MuI._2501_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6599_  (.A1(\MuI._0174_ ),
    .A2(\MuI._2500_ ),
    .B1(\MuI._2501_ ),
    .X(\MuI._2502_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6600_  (.A(\MuI._0141_ ),
    .B(\MuI._2502_ ),
    .X(\MuI._2503_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6601_  (.A(\MuI._2503_ ),
    .Y(\MuI._2504_ ));
 sky130_fd_sc_hd__nor3_4 \MuI._6602_  (.A(\MuI._0999_ ),
    .B(\MuI._2482_ ),
    .C(\MuI._2483_ ),
    .Y(\MuI._2505_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6603_  (.A_N(\MuI._1836_ ),
    .B(\MuI._1839_ ),
    .X(\MuI._2507_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6604_  (.A_N(\MuI._1839_ ),
    .B(\MuI._1836_ ),
    .X(\MuI._2508_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6605_  (.A(\MuI._2507_ ),
    .B(\MuI._2508_ ),
    .Y(\MuI._2509_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6606_  (.A_N(\MuI._1766_ ),
    .B(\MuI._1815_ ),
    .X(\MuI._2510_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6607_  (.A(\MuI._2510_ ),
    .Y(\MuI._2511_ ));
 sky130_fd_sc_hd__a22oi_1 \MuI._6608_  (.A1(\MuI._1795_ ),
    .A2(\MuI._1808_ ),
    .B1(\MuI._1831_ ),
    .B2(\MuI._2511_ ),
    .Y(\MuI._2512_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6609_  (.A(\MuI._1829_ ),
    .B(\MuI._2512_ ),
    .Y(\MuI._2513_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6610_  (.A1(\MuI._1814_ ),
    .A2(\MuI._2511_ ),
    .B1(\MuI._1809_ ),
    .Y(\MuI._2514_ ));
 sky130_fd_sc_hd__nor3b_1 \MuI._6611_  (.A(\MuI._1462_ ),
    .B(\MuI._1555_ ),
    .C_N(\MuI._1642_ ),
    .Y(\MuI._2515_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6612_  (.A1(\MuI._1642_ ),
    .A2(\MuI._1643_ ),
    .B1_N(\MuI._2515_ ),
    .X(\MuI._2516_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6613_  (.A0(\MuI._1645_ ),
    .A1(\MuI._2516_ ),
    .S(\MuI._1460_ ),
    .X(\MuI._2518_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6614_  (.A(\MuI._1290_ ),
    .B(\MuI._1457_ ),
    .X(\MuI._2519_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6615_  (.A(\MuI._1290_ ),
    .B(\MuI._1457_ ),
    .Y(\MuI._2520_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6616_  (.A(\MuI._1453_ ),
    .B_N(\MuI._1372_ ),
    .X(\MuI._2521_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6617_  (.A(\MuI._2521_ ),
    .B(\MuI._1452_ ),
    .Y(\MuI._2522_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6618_  (.A(\MuI._1447_ ),
    .B(\MuI._1449_ ),
    .X(\MuI._2523_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6619_  (.A(\MuI._1447_ ),
    .B(\MuI._1449_ ),
    .Y(\MuI._2524_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6620_  (.A(\MuI._2523_ ),
    .B(\MuI._2524_ ),
    .Y(\MuI._2525_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6621_  (.A(\MuI._1446_ ),
    .B_N(\MuI._1430_ ),
    .X(\MuI._2526_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6622_  (.A(\MuI._2526_ ),
    .B_N(\MuI._1445_ ),
    .X(\MuI._2527_ ));
 sky130_fd_sc_hd__nand4_1 \MuI._6623_  (.A(\MuI._2526_ ),
    .B(\MuI._1433_ ),
    .C(\MuI._1434_ ),
    .D(\MuI._1444_ ),
    .Y(\MuI._2529_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6624_  (.A1(\MuI._1436_ ),
    .A2(\MuI._1443_ ),
    .B1(\MuI._1426_ ),
    .Y(\MuI._2530_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6625_  (.A(\MuI._1413_ ),
    .B(\MuI._2530_ ),
    .Y(\MuI._2531_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6626_  (.A1(\MuI._3397_ ),
    .A2(\MuI._0421_ ),
    .B1(\MuI._1436_ ),
    .C1(\MuI._2531_ ),
    .X(\MuI._2532_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6627_  (.A1(\MuI._2527_ ),
    .A2(\MuI._2529_ ),
    .B1(\MuI._2532_ ),
    .X(\MuI._2533_ ));
 sky130_fd_sc_hd__a2111o_1 \MuI._6628_  (.A1(\MuI._2519_ ),
    .A2(\MuI._2520_ ),
    .B1(\MuI._2522_ ),
    .C1(\MuI._2525_ ),
    .D1(\MuI._2533_ ),
    .X(\MuI._2534_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6629_  (.A1(\MuI._1809_ ),
    .A2(\MuI._1814_ ),
    .B1(\MuI._1815_ ),
    .Y(\MuI._2535_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6630_  (.A(\MuI._1766_ ),
    .B(\MuI._2535_ ),
    .Y(\MuI._2536_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6631_  (.A1(\MuI._1460_ ),
    .A2(\MuI._1645_ ),
    .B1(\MuI._1764_ ),
    .X(\MuI._2537_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6632_  (.A(\MuI._1712_ ),
    .B(\MuI._2537_ ),
    .X(\MuI._2538_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6633_  (.A(\MuI._1712_ ),
    .B(\MuI._2537_ ),
    .Y(\MuI._2540_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._6634_  (.A1(\MuI._2511_ ),
    .A2(\MuI._2536_ ),
    .B1(\MuI._2538_ ),
    .B2(\MuI._2540_ ),
    .X(\MuI._2541_ ));
 sky130_fd_sc_hd__or4_1 \MuI._6635_  (.A(\MuI._2514_ ),
    .B(\MuI._2518_ ),
    .C(\MuI._2534_ ),
    .D(\MuI._2541_ ),
    .X(\MuI._2542_ ));
 sky130_fd_sc_hd__o21ai_1 \MuI._6636_  (.A1(\MuI._1712_ ),
    .A2(\MuI._2537_ ),
    .B1(\MuI._1762_ ),
    .Y(\MuI._2543_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6637_  (.A(\MuI._1760_ ),
    .B(\MuI._2543_ ),
    .Y(\MuI._2544_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6638_  (.A(\MuI._1438_ ),
    .B(\MuI._1442_ ),
    .Y(\MuI._2545_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6639_  (.A(\MuI._1454_ ),
    .B(\MuI._1456_ ),
    .Y(\MuI._2546_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6640_  (.A_N(\MuI._1238_ ),
    .B(\MuI._1458_ ),
    .X(\MuI._2547_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6641_  (.A(\MuI._2547_ ),
    .B(\MuI._1236_ ),
    .Y(\MuI._2548_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6642_  (.A(\MuI._1181_ ),
    .B(\MuI._2548_ ),
    .Y(\MuI._2549_ ));
 sky130_fd_sc_hd__o211ai_2 \MuI._6643_  (.A1(\MuI._1443_ ),
    .A2(\MuI._2545_ ),
    .B1(\MuI._2546_ ),
    .C1(\MuI._2549_ ),
    .Y(\MuI._2551_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6644_  (.A_N(\MuI._1458_ ),
    .B(\MuI._1238_ ),
    .X(\MuI._2552_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6645_  (.A(\MuI._2547_ ),
    .B(\MuI._2552_ ),
    .Y(\MuI._2553_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6646_  (.A(\MuI._1451_ ),
    .B_N(\MuI._1408_ ),
    .X(\MuI._2554_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6647_  (.A(\MuI._2554_ ),
    .B(\MuI._2523_ ),
    .Y(\MuI._2555_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6648_  (.A1(\MuI._3403_ ),
    .A2(\MuI._0421_ ),
    .B1(\MuI._1414_ ),
    .C1(\MuI._1441_ ),
    .X(\MuI._2556_ ));
 sky130_fd_sc_hd__or3_1 \MuI._6649_  (.A(\MuI._2553_ ),
    .B(\MuI._2555_ ),
    .C(\MuI._2556_ ),
    .X(\MuI._2557_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6650_  (.A(\MuI._2551_ ),
    .B(\MuI._2557_ ),
    .X(\MuI._2558_ ));
 sky130_fd_sc_hd__or4_4 \MuI._6651_  (.A(\MuI._2513_ ),
    .B(\MuI._2542_ ),
    .C(\MuI._2544_ ),
    .D(\MuI._2558_ ),
    .X(\MuI._2559_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6652_  (.A(\MuI._1829_ ),
    .B_N(\MuI._2512_ ),
    .X(\MuI._2560_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6653_  (.A1(\MuI._1827_ ),
    .A2(\MuI._1828_ ),
    .B1(\MuI._2560_ ),
    .X(\MuI._2562_ ));
 sky130_fd_sc_hd__xor2_4 \MuI._6654_  (.A(\MuI._1826_ ),
    .B(\MuI._2562_ ),
    .X(\MuI._2563_ ));
 sky130_fd_sc_hd__or3b_1 \MuI._6655_  (.A(\MuI._2553_ ),
    .B(\MuI._2555_ ),
    .C_N(\MuI._1442_ ),
    .X(\MuI._2564_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6656_  (.A1(\MuI._2557_ ),
    .A2(\MuI._2564_ ),
    .B1(\MuI._2544_ ),
    .C1(\MuI._2551_ ),
    .X(\MuI._2565_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6657_  (.A1(\MuI._2542_ ),
    .A2(\MuI._2565_ ),
    .B1(\MuI._2513_ ),
    .X(\MuI._2566_ ));
 sky130_fd_sc_hd__or4_1 \MuI._6658_  (.A(\MuI._0999_ ),
    .B(\MuI._2482_ ),
    .C(\MuI._2483_ ),
    .D(\MuI._2566_ ),
    .X(\MuI._2567_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._6659_  (.A1(\MuI._2505_ ),
    .A2(\MuI._2509_ ),
    .B1(\MuI._2559_ ),
    .C1(\MuI._2563_ ),
    .D1(\MuI._2567_ ),
    .X(\MuI._2568_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6660_  (.A(\MuI._0782_ ),
    .B(\MuI._2507_ ),
    .Y(\MuI._2569_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6661_  (.A(\MuI._1837_ ),
    .B(\MuI._2569_ ),
    .Y(\MuI._2570_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6662_  (.A0(\MuI._2509_ ),
    .A1(\MuI._2570_ ),
    .S(\MuI._2485_ ),
    .X(\MuI._2571_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6663_  (.A1(\MuI._1837_ ),
    .A2(\MuI._2507_ ),
    .B1(\MuI._0784_ ),
    .X(\MuI._2573_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6664_  (.A(\MuI._0550_ ),
    .B(\MuI._2573_ ),
    .X(\MuI._2574_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6665_  (.A0(\MuI._2570_ ),
    .A1(\MuI._2574_ ),
    .S(\MuI._2485_ ),
    .X(\MuI._2575_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6666_  (.A(\MuI._2568_ ),
    .B(\MuI._2571_ ),
    .C(\MuI._2575_ ),
    .X(\MuI._2576_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \MuI._6667_  (.A(\MuI._2576_ ),
    .X(\MuI._2577_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6668_  (.A1(\MuI._0550_ ),
    .A2(\MuI._2573_ ),
    .B1(\MuI._0547_ ),
    .Y(\MuI._2578_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6669_  (.A(\MuI._0549_ ),
    .B(\MuI._2578_ ),
    .Y(\MuI._2579_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6670_  (.A0(\MuI._2574_ ),
    .A1(\MuI._2579_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2580_ ));
 sky130_fd_sc_hd__o21ba_1 \MuI._6671_  (.A1(\MuI._1836_ ),
    .A2(\MuI._1840_ ),
    .B1_N(\MuI._0786_ ),
    .X(\MuI._2581_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6672_  (.A(\MuI._0282_ ),
    .B(\MuI._2581_ ),
    .Y(\MuI._2582_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6673_  (.A(\MuI._0282_ ),
    .B(\MuI._2581_ ),
    .Y(\MuI._2584_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6674_  (.A(\MuI._2582_ ),
    .B_N(\MuI._2584_ ),
    .X(\MuI._2585_ ));
 sky130_fd_sc_hd__clkinv_2 \MuI._6675_  (.A(\MuI._2585_ ),
    .Y(\MuI._2586_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6676_  (.A0(\MuI._2579_ ),
    .A1(\MuI._2586_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2587_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6677_  (.A(\MuI._2577_ ),
    .B(\MuI._2580_ ),
    .C(\MuI._2587_ ),
    .X(\MuI._2588_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6678_  (.A(\MuI._0787_ ),
    .B(\MuI._2582_ ),
    .Y(\MuI._2589_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6679_  (.A(\MuI._0147_ ),
    .B(\MuI._2589_ ),
    .Y(\MuI._2590_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6680_  (.A0(\MuI._2585_ ),
    .A1(\MuI._2590_ ),
    .S(\MuI._2485_ ),
    .X(\MuI._2591_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6681_  (.A1(\MuI._0146_ ),
    .A2(\MuI._0787_ ),
    .A3(\MuI._2582_ ),
    .B1(\MuI._0788_ ),
    .X(\MuI._2592_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6682_  (.A(\MuI._0013_ ),
    .B(\MuI._2592_ ),
    .Y(\MuI._2593_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6683_  (.A0(\MuI._2590_ ),
    .A1(\MuI._2593_ ),
    .S(\MuI._2485_ ),
    .X(\MuI._2595_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6684_  (.A(\MuI._2591_ ),
    .B(\MuI._2595_ ),
    .X(\MuI._2596_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6685_  (.A(\MuI._2596_ ),
    .Y(\MuI._2597_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6686_  (.A1(\MuI._0013_ ),
    .A2(\MuI._2592_ ),
    .B1_N(\MuI._0791_ ),
    .X(\MuI._2598_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6687_  (.A(\MuI._3304_ ),
    .B(\MuI._2598_ ),
    .Y(\MuI._2599_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6688_  (.A0(\MuI._2593_ ),
    .A1(\MuI._2599_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2600_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6689_  (.A(\MuI._2600_ ),
    .Y(\MuI._2601_ ));
 sky130_fd_sc_hd__a21boi_1 \MuI._6690_  (.A1(\MuI._0793_ ),
    .A2(\MuI._1841_ ),
    .B1_N(\MuI._2004_ ),
    .Y(\MuI._2602_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6691_  (.A1(\MuI._1996_ ),
    .A2(\MuI._2602_ ),
    .B1(\MuI._2394_ ),
    .Y(\MuI._2603_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6692_  (.A(\MuI._2383_ ),
    .B(\MuI._2603_ ),
    .X(\MuI._2604_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6693_  (.A(\MuI._2002_ ),
    .B(\MuI._2602_ ),
    .X(\MuI._2606_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6694_  (.A(\MuI._1996_ ),
    .B(\MuI._2606_ ),
    .Y(\MuI._2607_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6695_  (.A0(\MuI._2604_ ),
    .A1(\MuI._2607_ ),
    .S(\MuI._2505_ ),
    .X(\MuI._2608_ ));
 sky130_fd_sc_hd__and3b_1 \MuI._6696_  (.A_N(\MuI._2004_ ),
    .B(\MuI._0793_ ),
    .C(\MuI._1841_ ),
    .X(\MuI._2609_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6697_  (.A(\MuI._2602_ ),
    .B(\MuI._2609_ ),
    .X(\MuI._2610_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6698_  (.A1(\MuI._0999_ ),
    .A2(\MuI._2482_ ),
    .A3(\MuI._2483_ ),
    .B1(\MuI._2607_ ),
    .X(\MuI._2611_ ));
 sky130_fd_sc_hd__a211o_1 \MuI._6699_  (.A1(\MuI._2505_ ),
    .A2(\MuI._2599_ ),
    .B1(\MuI._2610_ ),
    .C1(\MuI._2611_ ),
    .X(\MuI._2612_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6700_  (.A_N(\MuI._2603_ ),
    .B(\MuI._2383_ ),
    .X(\MuI._2613_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6701_  (.A(\MuI._2391_ ),
    .B(\MuI._2613_ ),
    .Y(\MuI._2614_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6702_  (.A(\MuI._2380_ ),
    .B(\MuI._2614_ ),
    .X(\MuI._2615_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6703_  (.A0(\MuI._2604_ ),
    .A1(\MuI._2615_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2617_ ));
 sky130_fd_sc_hd__o21ai_2 \MuI._6704_  (.A1(\MuI._2384_ ),
    .A2(\MuI._2603_ ),
    .B1(\MuI._2392_ ),
    .Y(\MuI._2618_ ));
 sky130_fd_sc_hd__xor2_2 \MuI._6705_  (.A(\MuI._2366_ ),
    .B(\MuI._2618_ ),
    .X(\MuI._2619_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6706_  (.A0(\MuI._2615_ ),
    .A1(\MuI._2619_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2620_ ));
 sky130_fd_sc_hd__nor4_1 \MuI._6707_  (.A(\MuI._2608_ ),
    .B(\MuI._2612_ ),
    .C(\MuI._2617_ ),
    .D(\MuI._2620_ ),
    .Y(\MuI._2621_ ));
 sky130_fd_sc_hd__clkinv_2 \MuI._6708_  (.A(\MuI._2619_ ),
    .Y(\MuI._2622_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6709_  (.A(\MuI._2366_ ),
    .B_N(\MuI._2618_ ),
    .X(\MuI._2623_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6710_  (.A(\MuI._2364_ ),
    .B_N(\MuI._2623_ ),
    .X(\MuI._2624_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6711_  (.A(\MuI._2339_ ),
    .B(\MuI._2624_ ),
    .Y(\MuI._2625_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6712_  (.A0(\MuI._2622_ ),
    .A1(\MuI._2625_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2626_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6713_  (.A1(\MuI._2387_ ),
    .A2(\MuI._2623_ ),
    .B1(\MuI._2337_ ),
    .Y(\MuI._2628_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6714_  (.A(\MuI._2306_ ),
    .B(\MuI._2628_ ),
    .Y(\MuI._2629_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6715_  (.A0(\MuI._2625_ ),
    .A1(\MuI._2629_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2630_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6716_  (.A(\MuI._2621_ ),
    .B(\MuI._2626_ ),
    .C(\MuI._2630_ ),
    .X(\MuI._2631_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6717_  (.A(\MuI._2588_ ),
    .B(\MuI._2597_ ),
    .C(\MuI._2601_ ),
    .D(\MuI._2631_ ),
    .X(\MuI._2632_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6718_  (.A(\MuI._2306_ ),
    .B_N(\MuI._2628_ ),
    .X(\MuI._2633_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6719_  (.A(\MuI._2389_ ),
    .B(\MuI._2633_ ),
    .X(\MuI._2634_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6720_  (.A(\MuI._2241_ ),
    .B(\MuI._2634_ ),
    .X(\MuI._2635_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6721_  (.A0(\MuI._2629_ ),
    .A1(\MuI._2635_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2636_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6722_  (.A1(\MuI._2386_ ),
    .A2(\MuI._2398_ ),
    .B1(\MuI._2466_ ),
    .Y(\MuI._2637_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6723_  (.A(\MuI._2466_ ),
    .B(\MuI._2386_ ),
    .C(\MuI._2398_ ),
    .X(\MuI._2639_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6724_  (.A(\MuI._2637_ ),
    .B(\MuI._2639_ ),
    .Y(\MuI._2640_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6725_  (.A0(\MuI._2635_ ),
    .A1(\MuI._2640_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2641_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6726_  (.A(\MuI._2632_ ),
    .B(\MuI._2636_ ),
    .C(\MuI._2641_ ),
    .X(\MuI._2642_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._6727_  (.A(\MuI._2642_ ),
    .X(\MuI._2643_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6728_  (.A(\MuI._2464_ ),
    .B(\MuI._2637_ ),
    .X(\MuI._2644_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6729_  (.A(\MuI._2459_ ),
    .B(\MuI._2644_ ),
    .Y(\MuI._2645_ ));
 sky130_fd_sc_hd__clkinv_2 \MuI._6730_  (.A(\MuI._2645_ ),
    .Y(\MuI._2646_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6731_  (.A0(\MuI._2640_ ),
    .A1(\MuI._2646_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2647_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6732_  (.A1(\MuI._2637_ ),
    .A2(\MuI._2459_ ),
    .B1(\MuI._2469_ ),
    .Y(\MuI._2648_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6733_  (.A(\MuI._2444_ ),
    .B(\MuI._2648_ ),
    .Y(\MuI._2650_ ));
 sky130_fd_sc_hd__o21a_1 \MuI._6734_  (.A1(\MuI._2444_ ),
    .A2(\MuI._2648_ ),
    .B1(\MuI._2468_ ),
    .X(\MuI._2651_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6735_  (.A(\MuI._2424_ ),
    .B(\MuI._2651_ ),
    .Y(\MuI._2652_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6736_  (.A0(\MuI._2650_ ),
    .A1(\MuI._2652_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2653_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6737_  (.A0(\MuI._2645_ ),
    .A1(\MuI._2650_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2654_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6738_  (.A(\MuI._2653_ ),
    .B(\MuI._2654_ ),
    .Y(\MuI._2655_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6739_  (.A(\MuI._2643_ ),
    .B(\MuI._2647_ ),
    .C(\MuI._2655_ ),
    .X(\MuI._2656_ ));
 sky130_fd_sc_hd__clkinv_2 \MuI._6740_  (.A(\MuI._2652_ ),
    .Y(\MuI._2657_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6741_  (.A(\MuI._2474_ ),
    .B(\MuI._2467_ ),
    .C(\MuI._2471_ ),
    .X(\MuI._2658_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6742_  (.A(\MuI._2475_ ),
    .B(\MuI._2658_ ),
    .Y(\MuI._2659_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6743_  (.A0(\MuI._2657_ ),
    .A1(\MuI._2659_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2661_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6744_  (.A(\MuI._2308_ ),
    .B(\MuI._2475_ ),
    .Y(\MuI._2662_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6745_  (.A(\MuI._2476_ ),
    .B(\MuI._1747_ ),
    .Y(\MuI._2663_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6746_  (.A(\MuI._2662_ ),
    .B(\MuI._2663_ ),
    .Y(\MuI._2664_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6747_  (.A0(\MuI._2659_ ),
    .A1(\MuI._2664_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2665_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6748_  (.A(\MuI._2656_ ),
    .B(\MuI._2661_ ),
    .C(\MuI._2665_ ),
    .X(\MuI._2666_ ));
 sky130_fd_sc_hd__o31a_1 \MuI._6749_  (.A1(\MuI._1747_ ),
    .A2(\MuI._2308_ ),
    .A3(\MuI._2475_ ),
    .B1(\MuI._2477_ ),
    .X(\MuI._2667_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6750_  (.A(\MuI._2481_ ),
    .B(\MuI._2667_ ),
    .Y(\MuI._2668_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6751_  (.A(\MuI._2505_ ),
    .B(\MuI._2664_ ),
    .Y(\MuI._2669_ ));
 sky130_fd_sc_hd__o31ai_1 \MuI._6752_  (.A1(\MuI._2482_ ),
    .A2(\MuI._2505_ ),
    .A3(\MuI._2668_ ),
    .B1(\MuI._2669_ ),
    .Y(\MuI._2670_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6753_  (.A(\MuI._2666_ ),
    .B(\MuI._2670_ ),
    .Y(\MuI._2672_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6754_  (.A1(\MuI._2656_ ),
    .A2(\MuI._2661_ ),
    .B1(\MuI._2665_ ),
    .Y(\MuI._2673_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6755_  (.A(\MuI._2666_ ),
    .B(\MuI._2673_ ),
    .X(\MuI._2674_ ));
 sky130_fd_sc_hd__inv_2 \MuI._6756_  (.A(\MuI._2654_ ),
    .Y(\MuI._2675_ ));
 sky130_fd_sc_hd__nand3_1 \MuI._6757_  (.A(\MuI._2643_ ),
    .B(\MuI._2647_ ),
    .C(\MuI._2675_ ),
    .Y(\MuI._2676_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6758_  (.A1(\MuI._2643_ ),
    .A2(\MuI._2647_ ),
    .B1(\MuI._2675_ ),
    .X(\MuI._2677_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6759_  (.A(\MuI._2676_ ),
    .B(\MuI._2677_ ),
    .Y(\MuI._2678_ ));
 sky130_fd_sc_hd__and2_1 \MuI._6760_  (.A(\MuI._2621_ ),
    .B(\MuI._2626_ ),
    .X(\MuI._2679_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6761_  (.A(\MuI._2588_ ),
    .B(\MuI._2597_ ),
    .C(\MuI._2601_ ),
    .D(\MuI._2679_ ),
    .X(\MuI._2680_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6762_  (.A(\MuI._2588_ ),
    .B(\MuI._2597_ ),
    .C(\MuI._2601_ ),
    .X(\MuI._2681_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \MuI._6763_  (.A(\MuI._2681_ ),
    .X(\MuI._2683_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6764_  (.A1(\MuI._2683_ ),
    .A2(\MuI._2621_ ),
    .B1(\MuI._2626_ ),
    .Y(\MuI._2684_ ));
 sky130_fd_sc_hd__nand3_2 \MuI._6765_  (.A(\MuI._2577_ ),
    .B(\MuI._2580_ ),
    .C(\MuI._2587_ ),
    .Y(\MuI._2685_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6766_  (.A(\MuI._2608_ ),
    .B(\MuI._2612_ ),
    .X(\MuI._2686_ ));
 sky130_fd_sc_hd__or4_1 \MuI._6767_  (.A(\MuI._2685_ ),
    .B(\MuI._2596_ ),
    .C(\MuI._2600_ ),
    .D(\MuI._2686_ ),
    .X(\MuI._2687_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6768_  (.A(\MuI._2686_ ),
    .B(\MuI._2617_ ),
    .Y(\MuI._2688_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6769_  (.A(\MuI._2588_ ),
    .B(\MuI._2597_ ),
    .C(\MuI._2601_ ),
    .D(\MuI._2688_ ),
    .X(\MuI._2689_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6770_  (.A1(\MuI._2617_ ),
    .A2(\MuI._2687_ ),
    .B1(\MuI._2689_ ),
    .X(\MuI._2690_ ));
 sky130_fd_sc_hd__clkinv_2 \MuI._6771_  (.A(\MuI._2620_ ),
    .Y(\MuI._2691_ ));
 sky130_fd_sc_hd__a2bb2o_1 \MuI._6772_  (.A1_N(\MuI._2691_ ),
    .A2_N(\MuI._2689_ ),
    .B1(\MuI._2621_ ),
    .B2(\MuI._2683_ ),
    .X(\MuI._2692_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6773_  (.A(\MuI._2632_ ),
    .B(\MuI._2636_ ),
    .Y(\MuI._2694_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._6774_  (.A1(\MuI._2680_ ),
    .A2(\MuI._2684_ ),
    .B1(\MuI._2690_ ),
    .C1(\MuI._2692_ ),
    .D1(\MuI._2694_ ),
    .X(\MuI._2695_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6775_  (.A1(\MuI._2632_ ),
    .A2(\MuI._2636_ ),
    .B1(\MuI._2641_ ),
    .Y(\MuI._2696_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6776_  (.A0(\MuI._2599_ ),
    .A1(\MuI._2610_ ),
    .S(\MuI._2487_ ),
    .X(\MuI._2697_ ));
 sky130_fd_sc_hd__xor2_1 \MuI._6777_  (.A(\MuI._2683_ ),
    .B(\MuI._2697_ ),
    .X(\MuI._2698_ ));
 sky130_fd_sc_hd__or2_1 \MuI._6778_  (.A(\MuI._2685_ ),
    .B(\MuI._2591_ ),
    .X(\MuI._2699_ ));
 sky130_fd_sc_hd__a22o_1 \MuI._6779_  (.A1(\MuI._2588_ ),
    .A2(\MuI._2597_ ),
    .B1(\MuI._2699_ ),
    .B2(\MuI._2595_ ),
    .X(\MuI._2700_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6780_  (.A1(\MuI._2588_ ),
    .A2(\MuI._2597_ ),
    .B1(\MuI._2601_ ),
    .Y(\MuI._2701_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6781_  (.A(\MuI._2685_ ),
    .B(\MuI._2591_ ),
    .Y(\MuI._2702_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6782_  (.A1(\MuI._2577_ ),
    .A2(\MuI._2580_ ),
    .B1(\MuI._2587_ ),
    .X(\MuI._2703_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6783_  (.A(\MuI._2685_ ),
    .B(\MuI._2703_ ),
    .Y(\MuI._2705_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6784_  (.A1(\MuI._2568_ ),
    .A2(\MuI._2571_ ),
    .B1(\MuI._2575_ ),
    .Y(\MuI._2706_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6785_  (.A(\MuI._2577_ ),
    .B(\MuI._2706_ ),
    .Y(\MuI._2707_ ));
 sky130_fd_sc_hd__o211a_1 \MuI._6786_  (.A1(\MuI._2505_ ),
    .A2(\MuI._2563_ ),
    .B1(\MuI._2559_ ),
    .C1(\MuI._2567_ ),
    .X(\MuI._2708_ ));
 sky130_fd_sc_hd__mux2_1 \MuI._6787_  (.A0(\MuI._2563_ ),
    .A1(\MuI._2509_ ),
    .S(\MuI._2486_ ),
    .X(\MuI._2709_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6788_  (.A(\MuI._2708_ ),
    .B(\MuI._2709_ ),
    .Y(\MuI._2710_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6789_  (.A_N(\MuI.Exception ),
    .B(\MuI._2710_ ),
    .X(\MuI._2711_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6790_  (.A(\MuI._2568_ ),
    .B(\MuI._2571_ ),
    .Y(\MuI._2712_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6791_  (.A(\MuI._2577_ ),
    .B(\MuI._2580_ ),
    .Y(\MuI._2713_ ));
 sky130_fd_sc_hd__and4b_1 \MuI._6792_  (.A_N(\MuI._2707_ ),
    .B(\MuI._2711_ ),
    .C(\MuI._2712_ ),
    .D(\MuI._2713_ ),
    .X(\MuI._2714_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._6793_  (.A1(\MuI._2683_ ),
    .A2(\MuI._2701_ ),
    .B1(\MuI._2702_ ),
    .C1(\MuI._2705_ ),
    .D1(\MuI._2714_ ),
    .X(\MuI._2716_ ));
 sky130_fd_sc_hd__o2111a_1 \MuI._6794_  (.A1(\MuI._2643_ ),
    .A2(\MuI._2696_ ),
    .B1(\MuI._2698_ ),
    .C1(\MuI._2700_ ),
    .D1(\MuI._2716_ ),
    .X(\MuI._2717_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6795_  (.A(\MuI._2643_ ),
    .B(\MuI._2647_ ),
    .Y(\MuI._2718_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6796_  (.A1(\MuI._2505_ ),
    .A2(\MuI._2610_ ),
    .B1(\MuI._2611_ ),
    .X(\MuI._2719_ ));
 sky130_fd_sc_hd__or4_1 \MuI._6797_  (.A(\MuI._2685_ ),
    .B(\MuI._2596_ ),
    .C(\MuI._2600_ ),
    .D(\MuI._2697_ ),
    .X(\MuI._2720_ ));
 sky130_fd_sc_hd__or4_1 \MuI._6798_  (.A(\MuI._2685_ ),
    .B(\MuI._2596_ ),
    .C(\MuI._2600_ ),
    .D(\MuI._2612_ ),
    .X(\MuI._2721_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6799_  (.A1(\MuI._2719_ ),
    .A2(\MuI._2720_ ),
    .B1_N(\MuI._2721_ ),
    .X(\MuI._2722_ ));
 sky130_fd_sc_hd__o21bai_1 \MuI._6800_  (.A1(\MuI._2630_ ),
    .A2(\MuI._2680_ ),
    .B1_N(\MuI._2632_ ),
    .Y(\MuI._2723_ ));
 sky130_fd_sc_hd__a21bo_1 \MuI._6801_  (.A1(\MuI._2608_ ),
    .A2(\MuI._2721_ ),
    .B1_N(\MuI._2687_ ),
    .X(\MuI._2724_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6802_  (.A(\MuI._2722_ ),
    .B(\MuI._2723_ ),
    .C(\MuI._2724_ ),
    .X(\MuI._2725_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6803_  (.A(\MuI._2695_ ),
    .B(\MuI._2717_ ),
    .C(\MuI._2718_ ),
    .D(\MuI._2725_ ),
    .X(\MuI._2727_ ));
 sky130_fd_sc_hd__a21o_1 \MuI._6804_  (.A1(\MuI._2653_ ),
    .A2(\MuI._2676_ ),
    .B1(\MuI._2656_ ),
    .X(\MuI._2728_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6805_  (.A(\MuI._2656_ ),
    .B(\MuI._2661_ ),
    .Y(\MuI._2729_ ));
 sky130_fd_sc_hd__and4_1 \MuI._6806_  (.A(\MuI._2678_ ),
    .B(\MuI._2727_ ),
    .C(\MuI._2728_ ),
    .D(\MuI._2729_ ),
    .X(\MuI._2730_ ));
 sky130_fd_sc_hd__and3_1 \MuI._6807_  (.A(\MuI._2672_ ),
    .B(\MuI._2674_ ),
    .C(\MuI._2730_ ),
    .X(\MuI._2731_ ));
 sky130_fd_sc_hd__a21oi_2 \MuI._6808_  (.A1(\MuI._0141_ ),
    .A2(\MuI._2502_ ),
    .B1(\MuI._0130_ ),
    .Y(\MuI._2732_ ));
 sky130_fd_sc_hd__xor2_4 \MuI._6809_  (.A(\MuI._0086_ ),
    .B(\MuI._2732_ ),
    .X(\MuI._2733_ ));
 sky130_fd_sc_hd__or2b_1 \MuI._6810_  (.A(\MuI._2731_ ),
    .B_N(\MuI._2733_ ),
    .X(\MuI._2734_ ));
 sky130_fd_sc_hd__buf_2 \MuI._6811_  (.A(\MuI._2734_ ),
    .X(\MuI._2735_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6812_  (.A(\MuI._2504_ ),
    .B(\MuI._2735_ ),
    .Y(\MuI.Underflow ));
 sky130_fd_sc_hd__nor2_1 \MuI._6813_  (.A(\MuI._2503_ ),
    .B(\MuI._2735_ ),
    .Y(\MuI.Overflow ));
 sky130_fd_sc_hd__nor3_2 \MuI._6814_  (.A(\MuI.Exception ),
    .B(\MuI._2731_ ),
    .C(\MuI._2733_ ),
    .Y(\MuI._2737_ ));
 sky130_fd_sc_hd__clkbuf_2 \MuI._6815_  (.A(\MuI._2737_ ),
    .X(\MuI._2738_ ));
 sky130_fd_sc_hd__and2b_1 \MuI._6816_  (.A_N(\MuI._2710_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2739_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6817_  (.A(\MuI._2739_ ),
    .X(\MuI.result[0] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6818_  (.A_N(\MuI._2712_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2740_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6819_  (.A(\MuI._2740_ ),
    .X(\MuI.result[1] ));
 sky130_fd_sc_hd__and2_1 \MuI._6820_  (.A(\MuI._2707_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2741_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6821_  (.A(\MuI._2741_ ),
    .X(\MuI.result[2] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6822_  (.A_N(\MuI._2713_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2742_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6823_  (.A(\MuI._2742_ ),
    .X(\MuI.result[3] ));
 sky130_fd_sc_hd__and3_1 \MuI._6824_  (.A(\MuI._2685_ ),
    .B(\MuI._2703_ ),
    .C(\MuI._2737_ ),
    .X(\MuI._2744_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6825_  (.A(\MuI._2744_ ),
    .X(\MuI.result[4] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6826_  (.A_N(\MuI._2702_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2745_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6827_  (.A(\MuI._2745_ ),
    .X(\MuI.result[5] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6828_  (.A_N(\MuI._2700_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2746_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6829_  (.A(\MuI._2746_ ),
    .X(\MuI.result[6] ));
 sky130_fd_sc_hd__nor3b_1 \MuI._6830_  (.A(\MuI._2683_ ),
    .B(\MuI._2701_ ),
    .C_N(\MuI._2738_ ),
    .Y(\MuI.result[7] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6831_  (.A_N(\MuI._2698_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2747_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6832_  (.A(\MuI._2747_ ),
    .X(\MuI.result[8] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6833_  (.A_N(\MuI._2722_ ),
    .B(\MuI._2738_ ),
    .X(\MuI._2749_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6834_  (.A(\MuI._2749_ ),
    .X(\MuI.result[9] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6835_  (.A_N(\MuI._2724_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2750_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6836_  (.A(\MuI._2750_ ),
    .X(\MuI.result[10] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6837_  (.A_N(\MuI._2690_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2751_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6838_  (.A(\MuI._2751_ ),
    .X(\MuI.result[11] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6839_  (.A_N(\MuI._2692_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2752_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6840_  (.A(\MuI._2752_ ),
    .X(\MuI.result[12] ));
 sky130_fd_sc_hd__nor3b_1 \MuI._6841_  (.A(\MuI._2680_ ),
    .B(\MuI._2684_ ),
    .C_N(\MuI._2738_ ),
    .Y(\MuI.result[13] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6842_  (.A_N(\MuI._2723_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2753_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6843_  (.A(\MuI._2753_ ),
    .X(\MuI.result[14] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6844_  (.A_N(\MuI._2694_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2755_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6845_  (.A(\MuI._2755_ ),
    .X(\MuI.result[15] ));
 sky130_fd_sc_hd__or2_1 \MuI._6846_  (.A(\MuI.Exception ),
    .B(\MuI._2733_ ),
    .X(\MuI._2756_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \MuI._6847_  (.A(\MuI._2756_ ),
    .X(\MuI._2757_ ));
 sky130_fd_sc_hd__nor3_1 \MuI._6848_  (.A(\MuI._2643_ ),
    .B(\MuI._2696_ ),
    .C(\MuI._2757_ ),
    .Y(\MuI.result[16] ));
 sky130_fd_sc_hd__nor2_1 \MuI._6849_  (.A(\MuI._2718_ ),
    .B(\MuI._2757_ ),
    .Y(\MuI.result[17] ));
 sky130_fd_sc_hd__nor2_1 \MuI._6850_  (.A(\MuI._2678_ ),
    .B(\MuI._2757_ ),
    .Y(\MuI.result[18] ));
 sky130_fd_sc_hd__nor2_1 \MuI._6851_  (.A(\MuI._2728_ ),
    .B(\MuI._2757_ ),
    .Y(\MuI.result[19] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6852_  (.A_N(\MuI._2729_ ),
    .B(\MuI._2737_ ),
    .X(\MuI._2758_ ));
 sky130_fd_sc_hd__clkbuf_1 \MuI._6853_  (.A(\MuI._2758_ ),
    .X(\MuI.result[20] ));
 sky130_fd_sc_hd__nor2_1 \MuI._6854_  (.A(\MuI._2674_ ),
    .B(\MuI._2757_ ),
    .Y(\MuI.result[21] ));
 sky130_fd_sc_hd__nor2_1 \MuI._6855_  (.A(\MuI._2672_ ),
    .B(\MuI._2757_ ),
    .Y(\MuI.result[22] ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6856_  (.A(\MuI.b_operand[23] ),
    .B(\MuI._2489_ ),
    .Y(\MuI._2760_ ));
 sky130_fd_sc_hd__a211o_2 \MuI._6857_  (.A1(\MuI._2503_ ),
    .A2(\MuI._2733_ ),
    .B1(\MuI._2731_ ),
    .C1(\MuI.Exception ),
    .X(\MuI._2761_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6858_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2760_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[23] ));
 sky130_fd_sc_hd__or2b_1 \MuI._6859_  (.A(\MuI._2490_ ),
    .B_N(\MuI._2488_ ),
    .X(\MuI._2762_ ));
 sky130_fd_sc_hd__nand2_1 \MuI._6860_  (.A(\MuI.b_operand[23] ),
    .B(\MuI._2489_ ),
    .Y(\MuI._2763_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6861_  (.A(\MuI._2762_ ),
    .B(\MuI._2763_ ),
    .Y(\MuI._2764_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6862_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2764_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[24] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6863_  (.A_N(\MuI._2492_ ),
    .B(\MuI._0306_ ),
    .X(\MuI._2766_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6864_  (.A(\MuI._2766_ ),
    .B(\MuI._2491_ ),
    .Y(\MuI._2767_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6865_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2767_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[25] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6866_  (.A_N(\MuI._2494_ ),
    .B(\MuI._0273_ ),
    .X(\MuI._2768_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6867_  (.A(\MuI._2768_ ),
    .B(\MuI._2493_ ),
    .Y(\MuI._2769_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6868_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2769_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[26] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6869_  (.A_N(\MuI._2497_ ),
    .B(\MuI._0240_ ),
    .X(\MuI._2770_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6870_  (.A(\MuI._2770_ ),
    .B(\MuI._2496_ ),
    .Y(\MuI._2771_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6871_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2771_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[27] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6872_  (.A_N(\MuI._2499_ ),
    .B(\MuI._0207_ ),
    .X(\MuI._2772_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6873_  (.A(\MuI._2772_ ),
    .B(\MuI._2498_ ),
    .Y(\MuI._2774_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6874_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2774_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[28] ));
 sky130_fd_sc_hd__and2b_1 \MuI._6875_  (.A_N(\MuI._2501_ ),
    .B(\MuI._0174_ ),
    .X(\MuI._2775_ ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6876_  (.A(\MuI._2775_ ),
    .B(\MuI._2500_ ),
    .Y(\MuI._2776_ ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6877_  (.A1(\MuI._2735_ ),
    .A2(\MuI._2776_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[29] ));
 sky130_fd_sc_hd__a21oi_1 \MuI._6878_  (.A1(\MuI._2504_ ),
    .A2(\MuI._2735_ ),
    .B1(\MuI._2761_ ),
    .Y(\MuI.result[30] ));
 sky130_fd_sc_hd__xnor2_1 \MuI._6879_  (.A(\MuI.b_operand[31] ),
    .B(\MuI.a_operand[31] ),
    .Y(\MuI._2777_ ));
 sky130_fd_sc_hd__nor2_1 \MuI._6880_  (.A(\MuI.Exception ),
    .B(\MuI._2777_ ),
    .Y(\MuI.result[31] ));
 sky130_fd_sc_hd__buf_2 _06683_ (.A(net4),
    .X(_02020_));
 sky130_fd_sc_hd__nor2_2 _06684_ (.A(_02020_),
    .B(net3),
    .Y(_02031_));
 sky130_fd_sc_hd__buf_2 _06685_ (.A(_02031_),
    .X(_02042_));
 sky130_fd_sc_hd__buf_2 _06686_ (.A(_02042_),
    .X(_02053_));
 sky130_fd_sc_hd__buf_2 _06687_ (.A(net1),
    .X(_02064_));
 sky130_fd_sc_hd__nor2_2 _06688_ (.A(net2),
    .B(_02064_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_2 _06689_ (.A(_02053_),
    .B(_02075_),
    .Y(\AuI.AddBar_Sub ));
 sky130_fd_sc_hd__buf_4 _06690_ (.A(net37),
    .X(_02096_));
 sky130_fd_sc_hd__buf_4 _06691_ (.A(_02096_),
    .X(_02107_));
 sky130_fd_sc_hd__buf_6 _06692_ (.A(_02107_),
    .X(_02118_));
 sky130_fd_sc_hd__clkinv_2 _06693_ (.A(net2),
    .Y(_02129_));
 sky130_fd_sc_hd__and2_1 _06694_ (.A(_02129_),
    .B(net1),
    .X(_02140_));
 sky130_fd_sc_hd__buf_2 _06695_ (.A(_02140_),
    .X(_02151_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06696_ (.A(_02151_),
    .X(_02162_));
 sky130_fd_sc_hd__and3_1 _06697_ (.A(_02118_),
    .B(_02053_),
    .C(_02162_),
    .X(_02173_));
 sky130_fd_sc_hd__buf_2 _06698_ (.A(_02173_),
    .X(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__clkbuf_4 _06699_ (.A(net116),
    .X(_02194_));
 sky130_fd_sc_hd__buf_6 _06700_ (.A(_02194_),
    .X(_02205_));
 sky130_fd_sc_hd__clkbuf_8 _06701_ (.A(_02205_),
    .X(_02216_));
 sky130_fd_sc_hd__and3_1 _06702_ (.A(_02216_),
    .B(_02053_),
    .C(_02162_),
    .X(_02227_));
 sky130_fd_sc_hd__clkbuf_4 _06703_ (.A(_02227_),
    .X(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__buf_4 _06704_ (.A(net111),
    .X(_02248_));
 sky130_fd_sc_hd__clkbuf_8 _06705_ (.A(_02248_),
    .X(_02259_));
 sky130_fd_sc_hd__and3_1 _06706_ (.A(_02259_),
    .B(_02053_),
    .C(_02162_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_2 _06707_ (.A(_02270_),
    .X(\MuI.b_operand[2] ));
 sky130_fd_sc_hd__buf_4 _06708_ (.A(net110),
    .X(_02291_));
 sky130_fd_sc_hd__buf_4 _06709_ (.A(_02291_),
    .X(_02302_));
 sky130_fd_sc_hd__and3_1 _06710_ (.A(_02302_),
    .B(_02053_),
    .C(_02162_),
    .X(_02313_));
 sky130_fd_sc_hd__clkbuf_1 _06711_ (.A(_02313_),
    .X(\MuI.b_operand[3] ));
 sky130_fd_sc_hd__buf_2 _06712_ (.A(net109),
    .X(_02334_));
 sky130_fd_sc_hd__buf_4 _06713_ (.A(_02334_),
    .X(_02345_));
 sky130_fd_sc_hd__and3_1 _06714_ (.A(_02345_),
    .B(_02053_),
    .C(_02162_),
    .X(_02356_));
 sky130_fd_sc_hd__clkbuf_1 _06715_ (.A(_02356_),
    .X(\MuI.b_operand[4] ));
 sky130_fd_sc_hd__clkbuf_8 _06716_ (.A(net108),
    .X(_02377_));
 sky130_fd_sc_hd__buf_4 _06717_ (.A(_02377_),
    .X(_02388_));
 sky130_fd_sc_hd__and3_1 _06718_ (.A(_02388_),
    .B(_02053_),
    .C(_02162_),
    .X(_02399_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06719_ (.A(_02399_),
    .X(\MuI.b_operand[5] ));
 sky130_fd_sc_hd__clkbuf_8 _06720_ (.A(net107),
    .X(_02420_));
 sky130_fd_sc_hd__buf_4 _06721_ (.A(_02420_),
    .X(_02431_));
 sky130_fd_sc_hd__buf_4 _06722_ (.A(_02431_),
    .X(_02442_));
 sky130_fd_sc_hd__and3_1 _06723_ (.A(_02442_),
    .B(_02053_),
    .C(_02162_),
    .X(_02453_));
 sky130_fd_sc_hd__clkbuf_1 _06724_ (.A(_02453_),
    .X(\MuI.b_operand[6] ));
 sky130_fd_sc_hd__buf_4 _06725_ (.A(net66),
    .X(_02474_));
 sky130_fd_sc_hd__buf_4 _06726_ (.A(_02474_),
    .X(_02485_));
 sky130_fd_sc_hd__clkbuf_8 _06727_ (.A(_02485_),
    .X(_02496_));
 sky130_fd_sc_hd__and3_1 _06728_ (.A(_02496_),
    .B(_02053_),
    .C(_02162_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_1 _06729_ (.A(_02507_),
    .X(\MuI.b_operand[7] ));
 sky130_fd_sc_hd__buf_6 _06730_ (.A(net106),
    .X(_02528_));
 sky130_fd_sc_hd__buf_6 _06731_ (.A(_02528_),
    .X(_02539_));
 sky130_fd_sc_hd__buf_8 _06732_ (.A(_02539_),
    .X(_02550_));
 sky130_fd_sc_hd__and3_1 _06733_ (.A(_02550_),
    .B(_02053_),
    .C(_02162_),
    .X(_02561_));
 sky130_fd_sc_hd__clkbuf_2 _06734_ (.A(_02561_),
    .X(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__clkbuf_4 _06735_ (.A(net68),
    .X(_02582_));
 sky130_fd_sc_hd__buf_6 _06736_ (.A(_02582_),
    .X(_02593_));
 sky130_fd_sc_hd__buf_6 _06737_ (.A(_02593_),
    .X(_02604_));
 sky130_fd_sc_hd__clkbuf_2 _06738_ (.A(_02042_),
    .X(_02615_));
 sky130_fd_sc_hd__and3_1 _06739_ (.A(_02604_),
    .B(_02615_),
    .C(_02162_),
    .X(_02626_));
 sky130_fd_sc_hd__clkbuf_1 _06740_ (.A(_02626_),
    .X(\MuI.b_operand[9] ));
 sky130_fd_sc_hd__clkbuf_4 _06741_ (.A(net38),
    .X(_02647_));
 sky130_fd_sc_hd__buf_4 _06742_ (.A(_02647_),
    .X(_02658_));
 sky130_fd_sc_hd__buf_6 _06743_ (.A(_02658_),
    .X(_02669_));
 sky130_fd_sc_hd__clkbuf_2 _06744_ (.A(_02151_),
    .X(_02680_));
 sky130_fd_sc_hd__and3_1 _06745_ (.A(_02669_),
    .B(_02615_),
    .C(_02680_),
    .X(_02691_));
 sky130_fd_sc_hd__buf_2 _06746_ (.A(_02691_),
    .X(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__buf_6 _06747_ (.A(net39),
    .X(_02712_));
 sky130_fd_sc_hd__buf_6 _06748_ (.A(_02712_),
    .X(_02723_));
 sky130_fd_sc_hd__and3_1 _06749_ (.A(_02723_),
    .B(_02615_),
    .C(_02680_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_4 _06750_ (.A(_02734_),
    .X(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__buf_4 _06751_ (.A(net40),
    .X(_02754_));
 sky130_fd_sc_hd__buf_8 _06752_ (.A(_02754_),
    .X(_02765_));
 sky130_fd_sc_hd__and3_1 _06753_ (.A(_02765_),
    .B(_02615_),
    .C(_02680_),
    .X(_02776_));
 sky130_fd_sc_hd__clkbuf_1 _06754_ (.A(_02776_),
    .X(\MuI.b_operand[12] ));
 sky130_fd_sc_hd__buf_4 _06755_ (.A(net41),
    .X(_02797_));
 sky130_fd_sc_hd__buf_8 _06756_ (.A(_02797_),
    .X(_02808_));
 sky130_fd_sc_hd__and3_1 _06757_ (.A(_02808_),
    .B(_02615_),
    .C(_02680_),
    .X(_02819_));
 sky130_fd_sc_hd__clkbuf_1 _06758_ (.A(_02819_),
    .X(\MuI.b_operand[13] ));
 sky130_fd_sc_hd__buf_6 _06759_ (.A(net121),
    .X(_02840_));
 sky130_fd_sc_hd__buf_8 _06760_ (.A(_02840_),
    .X(_02851_));
 sky130_fd_sc_hd__buf_6 _06761_ (.A(_02851_),
    .X(_02862_));
 sky130_fd_sc_hd__and3_1 _06762_ (.A(_02862_),
    .B(_02615_),
    .C(_02680_),
    .X(_02873_));
 sky130_fd_sc_hd__clkbuf_4 _06763_ (.A(_02873_),
    .X(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__buf_4 _06764_ (.A(net43),
    .X(_02894_));
 sky130_fd_sc_hd__clkbuf_8 _06765_ (.A(_02894_),
    .X(_02905_));
 sky130_fd_sc_hd__buf_4 _06766_ (.A(_02905_),
    .X(_02916_));
 sky130_fd_sc_hd__and3_1 _06767_ (.A(_02916_),
    .B(_02615_),
    .C(_02680_),
    .X(_02927_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06768_ (.A(_02927_),
    .X(\MuI.b_operand[15] ));
 sky130_fd_sc_hd__clkbuf_4 _06769_ (.A(net44),
    .X(_02948_));
 sky130_fd_sc_hd__buf_6 _06770_ (.A(_02948_),
    .X(_02959_));
 sky130_fd_sc_hd__buf_6 _06771_ (.A(_02959_),
    .X(_02970_));
 sky130_fd_sc_hd__and3_1 _06772_ (.A(_02970_),
    .B(_02615_),
    .C(_02680_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _06773_ (.A(_02981_),
    .X(\MuI.b_operand[16] ));
 sky130_fd_sc_hd__buf_4 _06774_ (.A(net119),
    .X(_03002_));
 sky130_fd_sc_hd__buf_4 _06775_ (.A(_03002_),
    .X(_03013_));
 sky130_fd_sc_hd__buf_6 _06776_ (.A(_03013_),
    .X(_03024_));
 sky130_fd_sc_hd__and3_1 _06777_ (.A(_03024_),
    .B(_02615_),
    .C(_02680_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _06778_ (.A(_03035_),
    .X(\MuI.b_operand[17] ));
 sky130_fd_sc_hd__buf_4 _06779_ (.A(net118),
    .X(_03056_));
 sky130_fd_sc_hd__buf_6 _06780_ (.A(_03056_),
    .X(_03067_));
 sky130_fd_sc_hd__and3_1 _06781_ (.A(_03067_),
    .B(_02615_),
    .C(_02680_),
    .X(_03078_));
 sky130_fd_sc_hd__clkbuf_1 _06782_ (.A(_03078_),
    .X(\MuI.b_operand[18] ));
 sky130_fd_sc_hd__buf_4 _06783_ (.A(net117),
    .X(_03099_));
 sky130_fd_sc_hd__buf_6 _06784_ (.A(_03099_),
    .X(_03110_));
 sky130_fd_sc_hd__clkbuf_2 _06785_ (.A(_02042_),
    .X(_03121_));
 sky130_fd_sc_hd__and3_1 _06786_ (.A(_03110_),
    .B(_03121_),
    .C(_02680_),
    .X(_03131_));
 sky130_fd_sc_hd__clkbuf_2 _06787_ (.A(_03131_),
    .X(\MuI.b_operand[19] ));
 sky130_fd_sc_hd__buf_4 _06788_ (.A(net49),
    .X(_03152_));
 sky130_fd_sc_hd__clkbuf_8 _06789_ (.A(_03152_),
    .X(_03163_));
 sky130_fd_sc_hd__clkbuf_8 _06790_ (.A(_03163_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_2 _06791_ (.A(_02151_),
    .X(_03185_));
 sky130_fd_sc_hd__and3_1 _06792_ (.A(_03174_),
    .B(_03121_),
    .C(_03185_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_2 _06793_ (.A(_03196_),
    .X(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__buf_2 _06794_ (.A(net50),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_4 _06795_ (.A(_03217_),
    .X(_03228_));
 sky130_fd_sc_hd__clkbuf_8 _06796_ (.A(_03228_),
    .X(_03239_));
 sky130_fd_sc_hd__and3_1 _06797_ (.A(_03239_),
    .B(_03121_),
    .C(_03185_),
    .X(_03250_));
 sky130_fd_sc_hd__clkbuf_2 _06798_ (.A(_03250_),
    .X(\MuI.b_operand[21] ));
 sky130_fd_sc_hd__buf_2 _06799_ (.A(net51),
    .X(_03271_));
 sky130_fd_sc_hd__buf_4 _06800_ (.A(_03271_),
    .X(_03282_));
 sky130_fd_sc_hd__buf_4 _06801_ (.A(_03282_),
    .X(_03293_));
 sky130_fd_sc_hd__and3_1 _06802_ (.A(_03293_),
    .B(_03121_),
    .C(_03185_),
    .X(_03304_));
 sky130_fd_sc_hd__clkbuf_2 _06803_ (.A(_03304_),
    .X(\MuI.b_operand[22] ));
 sky130_fd_sc_hd__clkbuf_8 _06804_ (.A(net114),
    .X(_03324_));
 sky130_fd_sc_hd__buf_4 _06805_ (.A(_03324_),
    .X(_03335_));
 sky130_fd_sc_hd__buf_4 _06806_ (.A(_03335_),
    .X(_03346_));
 sky130_fd_sc_hd__and3_1 _06807_ (.A(_03346_),
    .B(_03121_),
    .C(_03185_),
    .X(_03357_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06808_ (.A(_03357_),
    .X(\MuI.b_operand[23] ));
 sky130_fd_sc_hd__buf_4 _06809_ (.A(net113),
    .X(_03378_));
 sky130_fd_sc_hd__buf_4 _06810_ (.A(_03378_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_4 _06811_ (.A(_03389_),
    .X(_03400_));
 sky130_fd_sc_hd__and3_1 _06812_ (.A(_03400_),
    .B(_03121_),
    .C(_03185_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _06813_ (.A(_03411_),
    .X(\MuI.b_operand[24] ));
 sky130_fd_sc_hd__clkbuf_4 _06814_ (.A(net54),
    .X(_03432_));
 sky130_fd_sc_hd__buf_4 _06815_ (.A(_03432_),
    .X(_03443_));
 sky130_fd_sc_hd__clkbuf_8 _06816_ (.A(_03443_),
    .X(_03454_));
 sky130_fd_sc_hd__and3_1 _06817_ (.A(_03454_),
    .B(_03121_),
    .C(_03185_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_1 _06818_ (.A(_03465_),
    .X(\MuI.b_operand[25] ));
 sky130_fd_sc_hd__buf_4 _06819_ (.A(net55),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_4 _06820_ (.A(_03486_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _06821_ (.A(_03497_),
    .X(_03507_));
 sky130_fd_sc_hd__and3_1 _06822_ (.A(_03507_),
    .B(_03121_),
    .C(_03185_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _06823_ (.A(_03518_),
    .X(\MuI.b_operand[26] ));
 sky130_fd_sc_hd__buf_2 _06824_ (.A(net112),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_4 _06825_ (.A(_03539_),
    .X(_03550_));
 sky130_fd_sc_hd__buf_4 _06826_ (.A(_03550_),
    .X(_03561_));
 sky130_fd_sc_hd__and3_1 _06827_ (.A(_03561_),
    .B(_03121_),
    .C(_03185_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _06828_ (.A(_03572_),
    .X(\MuI.b_operand[27] ));
 sky130_fd_sc_hd__buf_2 _06829_ (.A(net57),
    .X(_03593_));
 sky130_fd_sc_hd__buf_2 _06830_ (.A(_03593_),
    .X(_03604_));
 sky130_fd_sc_hd__clkbuf_4 _06831_ (.A(_03604_),
    .X(_03615_));
 sky130_fd_sc_hd__clkbuf_4 _06832_ (.A(_03615_),
    .X(_03626_));
 sky130_fd_sc_hd__and3_1 _06833_ (.A(_03626_),
    .B(_03121_),
    .C(_03185_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _06834_ (.A(_03637_),
    .X(\MuI.b_operand[28] ));
 sky130_fd_sc_hd__clkbuf_4 _06835_ (.A(net58),
    .X(_03658_));
 sky130_fd_sc_hd__clkbuf_4 _06836_ (.A(_03658_),
    .X(_03669_));
 sky130_fd_sc_hd__buf_2 _06837_ (.A(_03669_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_2 _06838_ (.A(_02042_),
    .X(_03690_));
 sky130_fd_sc_hd__and3_1 _06839_ (.A(_03680_),
    .B(_03690_),
    .C(_03185_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_1 _06840_ (.A(_03701_),
    .X(\MuI.b_operand[29] ));
 sky130_fd_sc_hd__buf_2 _06841_ (.A(net60),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_4 _06842_ (.A(_03722_),
    .X(_03733_));
 sky130_fd_sc_hd__clkbuf_4 _06843_ (.A(_03733_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_4 _06844_ (.A(_03744_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_2 _06845_ (.A(_02151_),
    .X(_03766_));
 sky130_fd_sc_hd__and3_1 _06846_ (.A(_03755_),
    .B(_03690_),
    .C(_03766_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_1 _06847_ (.A(_03777_),
    .X(\MuI.b_operand[30] ));
 sky130_fd_sc_hd__clkbuf_4 _06848_ (.A(net61),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_4 _06849_ (.A(_03798_),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_4 _06850_ (.A(_03809_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_4 _06851_ (.A(_03820_),
    .X(_03831_));
 sky130_fd_sc_hd__buf_4 _06852_ (.A(_03831_),
    .X(_03842_));
 sky130_fd_sc_hd__and3_1 _06853_ (.A(_03842_),
    .B(_03690_),
    .C(_03766_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _06854_ (.A(_03852_),
    .X(\MuI.b_operand[31] ));
 sky130_fd_sc_hd__clkbuf_4 _06855_ (.A(net115),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_4 _06856_ (.A(_03873_),
    .X(_03884_));
 sky130_fd_sc_hd__buf_4 _06857_ (.A(_03884_),
    .X(_03895_));
 sky130_fd_sc_hd__buf_4 _06858_ (.A(_03895_),
    .X(_03906_));
 sky130_fd_sc_hd__buf_4 _06859_ (.A(_03906_),
    .X(_03917_));
 sky130_fd_sc_hd__buf_4 _06860_ (.A(_03917_),
    .X(_03928_));
 sky130_fd_sc_hd__and3_1 _06861_ (.A(_03928_),
    .B(_03690_),
    .C(_03766_),
    .X(_03939_));
 sky130_fd_sc_hd__clkbuf_2 _06862_ (.A(_03939_),
    .X(\MuI.a_operand[0] ));
 sky130_fd_sc_hd__clkbuf_4 _06863_ (.A(net132),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_4 _06864_ (.A(_03960_),
    .X(_03971_));
 sky130_fd_sc_hd__buf_4 _06865_ (.A(_03971_),
    .X(_03982_));
 sky130_fd_sc_hd__clkbuf_4 _06866_ (.A(_03982_),
    .X(_03993_));
 sky130_fd_sc_hd__buf_4 _06867_ (.A(_03993_),
    .X(_04004_));
 sky130_fd_sc_hd__and3_1 _06868_ (.A(_04004_),
    .B(_03690_),
    .C(_03766_),
    .X(_04015_));
 sky130_fd_sc_hd__buf_2 _06869_ (.A(_04015_),
    .X(\MuI.a_operand[1] ));
 sky130_fd_sc_hd__clkbuf_4 _06870_ (.A(net127),
    .X(_04035_));
 sky130_fd_sc_hd__buf_4 _06871_ (.A(_04035_),
    .X(_04046_));
 sky130_fd_sc_hd__buf_6 _06872_ (.A(_04046_),
    .X(_04057_));
 sky130_fd_sc_hd__buf_4 _06873_ (.A(_04057_),
    .X(_04068_));
 sky130_fd_sc_hd__and3_1 _06874_ (.A(_04068_),
    .B(_03690_),
    .C(_03766_),
    .X(_04079_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06875_ (.A(_04079_),
    .X(\MuI.a_operand[2] ));
 sky130_fd_sc_hd__buf_2 _06876_ (.A(net126),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_4 _06877_ (.A(_04100_),
    .X(_04111_));
 sky130_fd_sc_hd__buf_4 _06878_ (.A(_04111_),
    .X(_04122_));
 sky130_fd_sc_hd__buf_4 _06879_ (.A(_04122_),
    .X(_04133_));
 sky130_fd_sc_hd__and3_1 _06880_ (.A(_04133_),
    .B(_03690_),
    .C(_03766_),
    .X(_04144_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06881_ (.A(_04144_),
    .X(\MuI.a_operand[3] ));
 sky130_fd_sc_hd__clkbuf_4 _06882_ (.A(net125),
    .X(_04165_));
 sky130_fd_sc_hd__buf_4 _06883_ (.A(_04165_),
    .X(_04176_));
 sky130_fd_sc_hd__buf_4 _06884_ (.A(_04176_),
    .X(_04186_));
 sky130_fd_sc_hd__buf_4 _06885_ (.A(_04186_),
    .X(_04197_));
 sky130_fd_sc_hd__and3_1 _06886_ (.A(_04197_),
    .B(_03690_),
    .C(_03766_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_2 _06887_ (.A(_04208_),
    .X(\MuI.a_operand[4] ));
 sky130_fd_sc_hd__clkbuf_4 _06888_ (.A(net124),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_4 _06889_ (.A(_04229_),
    .X(_04240_));
 sky130_fd_sc_hd__buf_4 _06890_ (.A(_04240_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_4 _06891_ (.A(_04251_),
    .X(_04262_));
 sky130_fd_sc_hd__and3_1 _06892_ (.A(_04262_),
    .B(_03690_),
    .C(_03766_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_2 _06893_ (.A(_04273_),
    .X(\MuI.a_operand[5] ));
 sky130_fd_sc_hd__buf_4 _06894_ (.A(net123),
    .X(_04294_));
 sky130_fd_sc_hd__buf_4 _06895_ (.A(_04294_),
    .X(_04305_));
 sky130_fd_sc_hd__buf_4 _06896_ (.A(_04305_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_4 _06897_ (.A(_04316_),
    .X(_04327_));
 sky130_fd_sc_hd__and3_1 _06898_ (.A(_04327_),
    .B(_03690_),
    .C(_03766_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_2 _06899_ (.A(_04338_),
    .X(\MuI.a_operand[6] ));
 sky130_fd_sc_hd__buf_4 _06900_ (.A(net34),
    .X(_04358_));
 sky130_fd_sc_hd__buf_4 _06901_ (.A(_04358_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_8 _06902_ (.A(_04369_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_4 _06903_ (.A(_04380_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_2 _06904_ (.A(_02031_),
    .X(_04402_));
 sky130_fd_sc_hd__and3_1 _06905_ (.A(_04391_),
    .B(_04402_),
    .C(_03766_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_2 _06906_ (.A(_04413_),
    .X(\MuI.a_operand[7] ));
 sky130_fd_sc_hd__buf_4 _06907_ (.A(net35),
    .X(_04434_));
 sky130_fd_sc_hd__buf_4 _06908_ (.A(_04434_),
    .X(_04445_));
 sky130_fd_sc_hd__buf_6 _06909_ (.A(_04445_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_4 _06910_ (.A(_04456_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_2 _06911_ (.A(_02151_),
    .X(_04478_));
 sky130_fd_sc_hd__and3_1 _06912_ (.A(_04467_),
    .B(_04402_),
    .C(_04478_),
    .X(_04489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06913_ (.A(_04489_),
    .X(\MuI.a_operand[8] ));
 sky130_fd_sc_hd__buf_4 _06914_ (.A(net36),
    .X(_04509_));
 sky130_fd_sc_hd__buf_6 _06915_ (.A(_04509_),
    .X(_04520_));
 sky130_fd_sc_hd__buf_6 _06916_ (.A(_04520_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_4 _06917_ (.A(_04531_),
    .X(_04542_));
 sky130_fd_sc_hd__and3_1 _06918_ (.A(_04542_),
    .B(_04402_),
    .C(_04478_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_2 _06919_ (.A(_04553_),
    .X(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__clkbuf_4 _06920_ (.A(net6),
    .X(_04574_));
 sky130_fd_sc_hd__buf_4 _06921_ (.A(_04574_),
    .X(_04585_));
 sky130_fd_sc_hd__buf_6 _06922_ (.A(_04585_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_4 _06923_ (.A(_04596_),
    .X(_04607_));
 sky130_fd_sc_hd__and3_1 _06924_ (.A(_04607_),
    .B(_04402_),
    .C(_04478_),
    .X(_04618_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06925_ (.A(_04618_),
    .X(\MuI.a_operand[10] ));
 sky130_fd_sc_hd__buf_4 _06926_ (.A(net7),
    .X(_04638_));
 sky130_fd_sc_hd__buf_4 _06927_ (.A(_04638_),
    .X(_04649_));
 sky130_fd_sc_hd__buf_4 _06928_ (.A(_04649_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_4 _06929_ (.A(_04660_),
    .X(_04671_));
 sky130_fd_sc_hd__and3_1 _06930_ (.A(_04671_),
    .B(_04402_),
    .C(_04478_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_2 _06931_ (.A(_04682_),
    .X(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__clkbuf_4 _06932_ (.A(net8),
    .X(_04703_));
 sky130_fd_sc_hd__buf_4 _06933_ (.A(_04703_),
    .X(_04714_));
 sky130_fd_sc_hd__buf_4 _06934_ (.A(_04714_),
    .X(_04725_));
 sky130_fd_sc_hd__buf_4 _06935_ (.A(_04725_),
    .X(_04736_));
 sky130_fd_sc_hd__and3_1 _06936_ (.A(_04736_),
    .B(_04402_),
    .C(_04478_),
    .X(_04747_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _06937_ (.A(_04747_),
    .X(\MuI.a_operand[12] ));
 sky130_fd_sc_hd__buf_2 _06938_ (.A(net9),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_8 _06939_ (.A(_04767_),
    .X(_04778_));
 sky130_fd_sc_hd__buf_6 _06940_ (.A(_04778_),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_4 _06941_ (.A(_04789_),
    .X(_04800_));
 sky130_fd_sc_hd__and3_1 _06942_ (.A(_04800_),
    .B(_04402_),
    .C(_04478_),
    .X(_04811_));
 sky130_fd_sc_hd__clkbuf_1 _06943_ (.A(_04811_),
    .X(\MuI.a_operand[13] ));
 sky130_fd_sc_hd__buf_4 _06944_ (.A(net10),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_8 _06945_ (.A(_04832_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_8 _06946_ (.A(_04843_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_4 _06947_ (.A(_04854_),
    .X(_04865_));
 sky130_fd_sc_hd__and3_1 _06948_ (.A(_04865_),
    .B(_04402_),
    .C(_04478_),
    .X(_04876_));
 sky130_fd_sc_hd__clkbuf_2 _06949_ (.A(_04876_),
    .X(\MuI.a_operand[14] ));
 sky130_fd_sc_hd__clkbuf_4 _06950_ (.A(net11),
    .X(_04896_));
 sky130_fd_sc_hd__buf_4 _06951_ (.A(_04896_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_8 _06952_ (.A(_04907_),
    .X(_04918_));
 sky130_fd_sc_hd__clkbuf_4 _06953_ (.A(_04918_),
    .X(_04929_));
 sky130_fd_sc_hd__and3_1 _06954_ (.A(_04929_),
    .B(_04402_),
    .C(_04478_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_2 _06955_ (.A(_04940_),
    .X(\MuI.a_operand[15] ));
 sky130_fd_sc_hd__buf_4 _06956_ (.A(net133),
    .X(_04961_));
 sky130_fd_sc_hd__buf_4 _06957_ (.A(_04961_),
    .X(_04972_));
 sky130_fd_sc_hd__buf_4 _06958_ (.A(_04972_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_4 _06959_ (.A(_04983_),
    .X(_04994_));
 sky130_fd_sc_hd__and3_1 _06960_ (.A(_04994_),
    .B(_04402_),
    .C(_04478_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_2 _06961_ (.A(_05005_),
    .X(\MuI.a_operand[16] ));
 sky130_fd_sc_hd__clkbuf_8 _06962_ (.A(net13),
    .X(_05025_));
 sky130_fd_sc_hd__buf_6 _06963_ (.A(_05025_),
    .X(_05036_));
 sky130_fd_sc_hd__buf_4 _06964_ (.A(_05036_),
    .X(_05047_));
 sky130_fd_sc_hd__clkbuf_4 _06965_ (.A(_05047_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_2 _06966_ (.A(_02031_),
    .X(_05069_));
 sky130_fd_sc_hd__and3_1 _06967_ (.A(_05058_),
    .B(_05069_),
    .C(_04478_),
    .X(_05080_));
 sky130_fd_sc_hd__buf_2 _06968_ (.A(_05080_),
    .X(\MuI.a_operand[17] ));
 sky130_fd_sc_hd__buf_4 _06969_ (.A(net14),
    .X(_05101_));
 sky130_fd_sc_hd__buf_4 _06970_ (.A(_05101_),
    .X(_05112_));
 sky130_fd_sc_hd__buf_4 _06971_ (.A(_05112_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_4 _06972_ (.A(_05123_),
    .X(_05134_));
 sky130_fd_sc_hd__clkbuf_2 _06973_ (.A(_02140_),
    .X(_05144_));
 sky130_fd_sc_hd__and3_1 _06974_ (.A(_05134_),
    .B(_05069_),
    .C(_05144_),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_2 _06975_ (.A(_05155_),
    .X(\MuI.a_operand[18] ));
 sky130_fd_sc_hd__clkbuf_4 _06976_ (.A(net15),
    .X(_05176_));
 sky130_fd_sc_hd__buf_4 _06977_ (.A(_05176_),
    .X(_05187_));
 sky130_fd_sc_hd__clkbuf_8 _06978_ (.A(_05187_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_4 _06979_ (.A(_05198_),
    .X(_05209_));
 sky130_fd_sc_hd__and3_1 _06980_ (.A(_05209_),
    .B(_05069_),
    .C(_05144_),
    .X(_05220_));
 sky130_fd_sc_hd__buf_2 _06981_ (.A(_05220_),
    .X(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__clkbuf_4 _06982_ (.A(net17),
    .X(_05241_));
 sky130_fd_sc_hd__buf_4 _06983_ (.A(_05241_),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_4 _06984_ (.A(_05252_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_4 _06985_ (.A(_05262_),
    .X(_05273_));
 sky130_fd_sc_hd__and3_1 _06986_ (.A(_05273_),
    .B(_05069_),
    .C(_05144_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_2 _06987_ (.A(_05284_),
    .X(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__clkbuf_4 _06988_ (.A(net18),
    .X(_05305_));
 sky130_fd_sc_hd__buf_4 _06989_ (.A(_05305_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_4 _06990_ (.A(_05316_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_4 _06991_ (.A(_05327_),
    .X(_05338_));
 sky130_fd_sc_hd__and3_1 _06992_ (.A(_05338_),
    .B(_05069_),
    .C(_05144_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _06993_ (.A(_05349_),
    .X(\MuI.a_operand[21] ));
 sky130_fd_sc_hd__clkbuf_4 _06994_ (.A(net19),
    .X(_05370_));
 sky130_fd_sc_hd__buf_4 _06995_ (.A(_05370_),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_4 _06996_ (.A(_05380_),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_4 _06997_ (.A(_05391_),
    .X(_05402_));
 sky130_fd_sc_hd__and3_1 _06998_ (.A(_05402_),
    .B(_05069_),
    .C(_05144_),
    .X(_05413_));
 sky130_fd_sc_hd__buf_2 _06999_ (.A(_05413_),
    .X(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__clkbuf_4 _07000_ (.A(net20),
    .X(_05434_));
 sky130_fd_sc_hd__buf_4 _07001_ (.A(_05434_),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_4 _07002_ (.A(_05445_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_4 _07003_ (.A(_05456_),
    .X(_05467_));
 sky130_fd_sc_hd__and3_1 _07004_ (.A(_05467_),
    .B(_05069_),
    .C(_05144_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_2 _07005_ (.A(_05478_),
    .X(\MuI.a_operand[23] ));
 sky130_fd_sc_hd__clkbuf_4 _07006_ (.A(net21),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_4 _07007_ (.A(_05498_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_4 _07008_ (.A(_05509_),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_4 _07009_ (.A(_05520_),
    .X(_05531_));
 sky130_fd_sc_hd__and3_1 _07010_ (.A(_05531_),
    .B(_05069_),
    .C(_05144_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_2 _07011_ (.A(_05542_),
    .X(\MuI.a_operand[24] ));
 sky130_fd_sc_hd__clkbuf_4 _07012_ (.A(net22),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_4 _07013_ (.A(_05563_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_4 _07014_ (.A(_05574_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_4 _07015_ (.A(_05585_),
    .X(_05595_));
 sky130_fd_sc_hd__and3_1 _07016_ (.A(_05595_),
    .B(_05069_),
    .C(_05144_),
    .X(_05606_));
 sky130_fd_sc_hd__buf_4 _07017_ (.A(_05606_),
    .X(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__clkbuf_4 _07018_ (.A(net23),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_4 _07019_ (.A(_05627_),
    .X(_05638_));
 sky130_fd_sc_hd__buf_4 _07020_ (.A(_05638_),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_4 _07021_ (.A(_05649_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_4 _07022_ (.A(_05660_),
    .X(_05671_));
 sky130_fd_sc_hd__and3_1 _07023_ (.A(_05671_),
    .B(_05069_),
    .C(_05144_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_2 _07024_ (.A(_05682_),
    .X(\MuI.a_operand[26] ));
 sky130_fd_sc_hd__buf_4 _07025_ (.A(net130),
    .X(_05702_));
 sky130_fd_sc_hd__buf_2 _07026_ (.A(_05702_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_4 _07027_ (.A(_05713_),
    .X(_05724_));
 sky130_fd_sc_hd__and3_1 _07028_ (.A(_05724_),
    .B(_02042_),
    .C(_05144_),
    .X(_05735_));
 sky130_fd_sc_hd__clkbuf_2 _07029_ (.A(_05735_),
    .X(\MuI.a_operand[27] ));
 sky130_fd_sc_hd__clkbuf_4 _07030_ (.A(net25),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_4 _07031_ (.A(_05756_),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_4 _07032_ (.A(_05767_),
    .X(_05777_));
 sky130_fd_sc_hd__clkbuf_4 _07033_ (.A(_05777_),
    .X(_05788_));
 sky130_fd_sc_hd__and3_1 _07034_ (.A(_05788_),
    .B(_02042_),
    .C(_02151_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_2 _07035_ (.A(_05799_),
    .X(\MuI.a_operand[28] ));
 sky130_fd_sc_hd__clkbuf_4 _07036_ (.A(net128),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_4 _07037_ (.A(_05820_),
    .X(_05831_));
 sky130_fd_sc_hd__clkbuf_4 _07038_ (.A(_05831_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_4 _07039_ (.A(_05842_),
    .X(_05853_));
 sky130_fd_sc_hd__and3_1 _07040_ (.A(_05853_),
    .B(_02042_),
    .C(_02151_),
    .X(_05863_));
 sky130_fd_sc_hd__clkbuf_2 _07041_ (.A(_05863_),
    .X(\MuI.a_operand[29] ));
 sky130_fd_sc_hd__clkbuf_4 _07042_ (.A(net28),
    .X(_05884_));
 sky130_fd_sc_hd__buf_4 _07043_ (.A(_05884_),
    .X(_05895_));
 sky130_fd_sc_hd__clkbuf_4 _07044_ (.A(_05895_),
    .X(_05906_));
 sky130_fd_sc_hd__clkbuf_4 _07045_ (.A(_05906_),
    .X(_05917_));
 sky130_fd_sc_hd__and3_1 _07046_ (.A(_05917_),
    .B(_02042_),
    .C(_02151_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_2 _07047_ (.A(_05928_),
    .X(\MuI.a_operand[30] ));
 sky130_fd_sc_hd__clkbuf_4 _07048_ (.A(net29),
    .X(_05948_));
 sky130_fd_sc_hd__buf_4 _07049_ (.A(_05948_),
    .X(_05959_));
 sky130_fd_sc_hd__buf_4 _07050_ (.A(_05959_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_4 _07051_ (.A(_05970_),
    .X(_05981_));
 sky130_fd_sc_hd__buf_2 _07052_ (.A(_05981_),
    .X(_05992_));
 sky130_fd_sc_hd__and3_1 _07053_ (.A(_05992_),
    .B(_02042_),
    .C(_02151_),
    .X(_06003_));
 sky130_fd_sc_hd__clkbuf_1 _07054_ (.A(_06003_),
    .X(\MuI.a_operand[31] ));
 sky130_fd_sc_hd__buf_2 _07055_ (.A(net3),
    .X(_06023_));
 sky130_fd_sc_hd__and3b_1 _07056_ (.A_N(_06023_),
    .B(_02140_),
    .C(_02020_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_4 _07057_ (.A(_06034_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_4 _07058_ (.A(_06045_),
    .X(_06056_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07059_ (.A(_06056_),
    .X(_06067_));
 sky130_fd_sc_hd__and2_1 _07062_ (.A(_04004_),
    .B(_06067_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _07063_ (.A(_06098_),
    .X(\FuI.a_operand[1] ));
 sky130_fd_sc_hd__and2_1 _07064_ (.A(_04068_),
    .B(_06067_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_1 _07065_ (.A(_06119_),
    .X(\FuI.a_operand[2] ));
 sky130_fd_sc_hd__and2_1 _07066_ (.A(_04133_),
    .B(_06067_),
    .X(_06140_));
 sky130_fd_sc_hd__clkbuf_1 _07067_ (.A(_06140_),
    .X(\FuI.a_operand[3] ));
 sky130_fd_sc_hd__and2_1 _07068_ (.A(_04197_),
    .B(_06067_),
    .X(_06160_));
 sky130_fd_sc_hd__clkbuf_1 _07069_ (.A(_06160_),
    .X(\FuI.a_operand[4] ));
 sky130_fd_sc_hd__and2_1 _07070_ (.A(_04262_),
    .B(_06067_),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _07071_ (.A(_06181_),
    .X(\FuI.a_operand[5] ));
 sky130_fd_sc_hd__and2_1 _07072_ (.A(_04327_),
    .B(_06067_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _07073_ (.A(_06202_),
    .X(\FuI.a_operand[6] ));
 sky130_fd_sc_hd__and2_1 _07074_ (.A(_04391_),
    .B(_06067_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _07075_ (.A(_06222_),
    .X(\FuI.a_operand[7] ));
 sky130_fd_sc_hd__and2_1 _07076_ (.A(_04467_),
    .B(_06067_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _07077_ (.A(_06243_),
    .X(\FuI.a_operand[8] ));
 sky130_fd_sc_hd__and2_1 _07078_ (.A(_04542_),
    .B(_06067_),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _07079_ (.A(_06264_),
    .X(\FuI.a_operand[9] ));
 sky130_fd_sc_hd__clkbuf_2 _07080_ (.A(_06056_),
    .X(_06284_));
 sky130_fd_sc_hd__and2_1 _07081_ (.A(_04607_),
    .B(_06284_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_1 _07082_ (.A(_06295_),
    .X(\FuI.a_operand[10] ));
 sky130_fd_sc_hd__and2_1 _07083_ (.A(_04671_),
    .B(_06284_),
    .X(_06316_));
 sky130_fd_sc_hd__clkbuf_1 _07084_ (.A(_06316_),
    .X(\FuI.a_operand[11] ));
 sky130_fd_sc_hd__and2_1 _07085_ (.A(_04736_),
    .B(_06284_),
    .X(_06336_));
 sky130_fd_sc_hd__clkbuf_1 _07086_ (.A(_06336_),
    .X(\FuI.a_operand[12] ));
 sky130_fd_sc_hd__and2_1 _07087_ (.A(_04800_),
    .B(_06284_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _07088_ (.A(_06356_),
    .X(\FuI.a_operand[13] ));
 sky130_fd_sc_hd__and2_1 _07089_ (.A(_04865_),
    .B(_06284_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _07090_ (.A(_06377_),
    .X(\FuI.a_operand[14] ));
 sky130_fd_sc_hd__and2_1 _07091_ (.A(_04929_),
    .B(_06284_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _07092_ (.A(_06397_),
    .X(\FuI.a_operand[15] ));
 sky130_fd_sc_hd__and2_1 _07093_ (.A(_04994_),
    .B(_06284_),
    .X(_06410_));
 sky130_fd_sc_hd__clkbuf_1 _07094_ (.A(_06410_),
    .X(\FuI.a_operand[16] ));
 sky130_fd_sc_hd__and2_1 _07095_ (.A(_05058_),
    .B(_06284_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _07096_ (.A(_06411_),
    .X(\FuI.a_operand[17] ));
 sky130_fd_sc_hd__and2_1 _07097_ (.A(_05134_),
    .B(_06284_),
    .X(_06412_));
 sky130_fd_sc_hd__clkbuf_1 _07098_ (.A(_06412_),
    .X(\FuI.a_operand[18] ));
 sky130_fd_sc_hd__and2_1 _07099_ (.A(_05209_),
    .B(_06284_),
    .X(_06413_));
 sky130_fd_sc_hd__clkbuf_1 _07100_ (.A(_06413_),
    .X(\FuI.a_operand[19] ));
 sky130_fd_sc_hd__clkbuf_2 _07101_ (.A(_06056_),
    .X(_06414_));
 sky130_fd_sc_hd__and2_1 _07102_ (.A(_05273_),
    .B(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _07103_ (.A(_06415_),
    .X(\FuI.a_operand[20] ));
 sky130_fd_sc_hd__and2_1 _07104_ (.A(_05338_),
    .B(_06414_),
    .X(_06416_));
 sky130_fd_sc_hd__clkbuf_1 _07105_ (.A(_06416_),
    .X(\FuI.a_operand[21] ));
 sky130_fd_sc_hd__and2_1 _07106_ (.A(_05402_),
    .B(_06414_),
    .X(_06417_));
 sky130_fd_sc_hd__clkbuf_1 _07107_ (.A(_06417_),
    .X(\FuI.a_operand[22] ));
 sky130_fd_sc_hd__and2_1 _07108_ (.A(_05467_),
    .B(_06414_),
    .X(_06418_));
 sky130_fd_sc_hd__clkbuf_2 _07109_ (.A(_06418_),
    .X(\FuI.a_operand[23] ));
 sky130_fd_sc_hd__and2_1 _07110_ (.A(_05531_),
    .B(_06414_),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_1 _07111_ (.A(_06419_),
    .X(\FuI.a_operand[24] ));
 sky130_fd_sc_hd__and2_1 _07112_ (.A(_05595_),
    .B(_06414_),
    .X(_06420_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07113_ (.A(_06420_),
    .X(\FuI.a_operand[25] ));
 sky130_fd_sc_hd__and2_1 _07114_ (.A(_05671_),
    .B(_06414_),
    .X(_06421_));
 sky130_fd_sc_hd__clkbuf_2 _07115_ (.A(_06421_),
    .X(\FuI.a_operand[26] ));
 sky130_fd_sc_hd__and2_1 _07116_ (.A(_05724_),
    .B(_06414_),
    .X(_06422_));
 sky130_fd_sc_hd__clkbuf_1 _07117_ (.A(_06422_),
    .X(\FuI.a_operand[27] ));
 sky130_fd_sc_hd__and2_1 _07118_ (.A(_05788_),
    .B(_06414_),
    .X(_06423_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07119_ (.A(_06423_),
    .X(\FuI.a_operand[28] ));
 sky130_fd_sc_hd__and2_1 _07120_ (.A(_05853_),
    .B(_06414_),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _07121_ (.A(_06424_),
    .X(\FuI.a_operand[29] ));
 sky130_fd_sc_hd__and2_1 _07122_ (.A(_05917_),
    .B(_06056_),
    .X(_06425_));
 sky130_fd_sc_hd__clkbuf_1 _07123_ (.A(_06425_),
    .X(\FuI.a_operand[30] ));
 sky130_fd_sc_hd__and2_1 _07124_ (.A(_05992_),
    .B(_06056_),
    .X(_06426_));
 sky130_fd_sc_hd__clkbuf_1 _07125_ (.A(_06426_),
    .X(\FuI.a_operand[31] ));
 sky130_fd_sc_hd__nand3_2 _07126_ (.A(_02020_),
    .B(_06023_),
    .C(_02140_),
    .Y(_06427_));
 sky130_fd_sc_hd__clkbuf_8 _07127_ (.A(_06427_),
    .X(_06428_));
 sky130_fd_sc_hd__clkbuf_4 _07128_ (.A(net60),
    .X(_06429_));
 sky130_fd_sc_hd__buf_2 _07129_ (.A(net127),
    .X(_06430_));
 sky130_fd_sc_hd__clkbuf_4 _07130_ (.A(net126),
    .X(_06431_));
 sky130_fd_sc_hd__and4_1 _07131_ (.A(net112),
    .B(_03593_),
    .C(_06430_),
    .D(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_4 _07132_ (.A(_04100_),
    .X(_06433_));
 sky130_fd_sc_hd__buf_2 _07133_ (.A(net112),
    .X(_06434_));
 sky130_fd_sc_hd__a22oi_1 _07134_ (.A1(_03604_),
    .A2(_04035_),
    .B1(_06433_),
    .B2(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__buf_4 _07135_ (.A(net132),
    .X(_06436_));
 sky130_fd_sc_hd__buf_4 _07136_ (.A(_06436_),
    .X(_06437_));
 sky130_fd_sc_hd__and4bb_1 _07137_ (.A_N(_06432_),
    .B_N(_06435_),
    .C(net58),
    .D(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__buf_2 _07138_ (.A(net58),
    .X(_06439_));
 sky130_fd_sc_hd__o2bb2a_1 _07139_ (.A1_N(_06439_),
    .A2_N(_06437_),
    .B1(_06432_),
    .B2(_06435_),
    .X(_06440_));
 sky130_fd_sc_hd__nor2_1 _07140_ (.A(_06438_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__clkbuf_4 _07141_ (.A(_03593_),
    .X(_06442_));
 sky130_fd_sc_hd__buf_4 _07142_ (.A(_04035_),
    .X(_06443_));
 sky130_fd_sc_hd__buf_2 _07143_ (.A(net112),
    .X(_06444_));
 sky130_fd_sc_hd__a22o_1 _07144_ (.A1(_06442_),
    .A2(_03960_),
    .B1(_06443_),
    .B2(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__buf_4 _07145_ (.A(net127),
    .X(_06446_));
 sky130_fd_sc_hd__and4_1 _07146_ (.A(_06444_),
    .B(_06442_),
    .C(_03960_),
    .D(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__a31o_1 _07147_ (.A1(_03658_),
    .A2(_03873_),
    .A3(_06445_),
    .B1(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__xor2_1 _07148_ (.A(_06441_),
    .B(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__and3_1 _07149_ (.A(_06429_),
    .B(_03906_),
    .C(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__a21oi_1 _07150_ (.A1(_03733_),
    .A2(_03906_),
    .B1(_06449_),
    .Y(_06451_));
 sky130_fd_sc_hd__nor2_2 _07151_ (.A(_06450_),
    .B(_06451_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _07152_ (.A(_03669_),
    .B(_03895_),
    .Y(_06453_));
 sky130_fd_sc_hd__and2b_1 _07153_ (.A_N(_06447_),
    .B(_06445_),
    .X(_06454_));
 sky130_fd_sc_hd__xnor2_2 _07154_ (.A(_06453_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__and4_2 _07155_ (.A(_03561_),
    .B(_03615_),
    .C(_03895_),
    .D(_03993_),
    .X(_06456_));
 sky130_fd_sc_hd__and2_1 _07156_ (.A(_06455_),
    .B(_06456_),
    .X(_06457_));
 sky130_fd_sc_hd__and2_1 _07157_ (.A(_06452_),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__and4_1 _07158_ (.A(_02096_),
    .B(_02194_),
    .C(net23),
    .D(net130),
    .X(_06459_));
 sky130_fd_sc_hd__buf_4 _07159_ (.A(net111),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_4 _07160_ (.A(net22),
    .X(_06461_));
 sky130_fd_sc_hd__nand2_1 _07161_ (.A(_06460_),
    .B(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__buf_6 _07162_ (.A(net116),
    .X(_06463_));
 sky130_fd_sc_hd__a22oi_2 _07163_ (.A1(_06463_),
    .A2(_05627_),
    .B1(net130),
    .B2(_02107_),
    .Y(_06464_));
 sky130_fd_sc_hd__or3_1 _07164_ (.A(_06459_),
    .B(_06462_),
    .C(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__buf_2 _07165_ (.A(net21),
    .X(_06466_));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(_06460_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__a22oi_2 _07167_ (.A1(_06463_),
    .A2(_06461_),
    .B1(_05627_),
    .B2(_02107_),
    .Y(_06468_));
 sky130_fd_sc_hd__buf_4 _07168_ (.A(net37),
    .X(_06469_));
 sky130_fd_sc_hd__and4_1 _07169_ (.A(_06469_),
    .B(_02194_),
    .C(net22),
    .D(_05627_),
    .X(_06470_));
 sky130_fd_sc_hd__o21bai_1 _07170_ (.A1(_06467_),
    .A2(_06468_),
    .B1_N(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__o21ai_1 _07171_ (.A1(_06459_),
    .A2(_06464_),
    .B1(_06462_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand3_1 _07172_ (.A(_06465_),
    .B(_06471_),
    .C(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__a21o_1 _07173_ (.A1(_06465_),
    .A2(_06472_),
    .B1(_06471_),
    .X(_06474_));
 sky130_fd_sc_hd__clkbuf_8 _07174_ (.A(net108),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_4 _07175_ (.A(net19),
    .X(_06476_));
 sky130_fd_sc_hd__buf_4 _07176_ (.A(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__nand2_1 _07177_ (.A(_06475_),
    .B(_06477_),
    .Y(_06478_));
 sky130_fd_sc_hd__buf_4 _07178_ (.A(net110),
    .X(_06479_));
 sky130_fd_sc_hd__buf_4 _07179_ (.A(net109),
    .X(_06480_));
 sky130_fd_sc_hd__and4_1 _07180_ (.A(_06479_),
    .B(_06480_),
    .C(net20),
    .D(_06466_),
    .X(_06481_));
 sky130_fd_sc_hd__a22o_1 _07181_ (.A1(_06480_),
    .A2(_05434_),
    .B1(_06466_),
    .B2(_06479_),
    .X(_06482_));
 sky130_fd_sc_hd__and2b_1 _07182_ (.A_N(_06481_),
    .B(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__xnor2_1 _07183_ (.A(_06478_),
    .B(_06483_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand3_1 _07184_ (.A(_06473_),
    .B(_06474_),
    .C(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__or3_1 _07185_ (.A(_06470_),
    .B(_06467_),
    .C(_06468_),
    .X(_06486_));
 sky130_fd_sc_hd__o21ai_1 _07186_ (.A1(_06470_),
    .A2(_06468_),
    .B1(_06467_),
    .Y(_06487_));
 sky130_fd_sc_hd__buf_4 _07187_ (.A(net111),
    .X(_06488_));
 sky130_fd_sc_hd__clkbuf_4 _07188_ (.A(net20),
    .X(_06489_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_06488_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__buf_6 _07190_ (.A(net116),
    .X(_06491_));
 sky130_fd_sc_hd__buf_6 _07191_ (.A(_02096_),
    .X(_06492_));
 sky130_fd_sc_hd__a22oi_2 _07192_ (.A1(_06491_),
    .A2(_06466_),
    .B1(_06461_),
    .B2(_06492_),
    .Y(_06493_));
 sky130_fd_sc_hd__buf_4 _07193_ (.A(net37),
    .X(_06494_));
 sky130_fd_sc_hd__buf_4 _07194_ (.A(net116),
    .X(_06495_));
 sky130_fd_sc_hd__and4_1 _07195_ (.A(_06494_),
    .B(_06495_),
    .C(net21),
    .D(_06461_),
    .X(_06496_));
 sky130_fd_sc_hd__o21bai_1 _07196_ (.A1(_06490_),
    .A2(_06493_),
    .B1_N(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__a21o_1 _07197_ (.A1(_06486_),
    .A2(_06487_),
    .B1(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__nand2_1 _07198_ (.A(_06475_),
    .B(_05316_),
    .Y(_06499_));
 sky130_fd_sc_hd__buf_4 _07199_ (.A(net109),
    .X(_06500_));
 sky130_fd_sc_hd__buf_4 _07200_ (.A(net110),
    .X(_06501_));
 sky130_fd_sc_hd__a22oi_1 _07201_ (.A1(_06500_),
    .A2(_06476_),
    .B1(_06489_),
    .B2(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__buf_4 _07202_ (.A(net110),
    .X(_06503_));
 sky130_fd_sc_hd__buf_4 _07203_ (.A(net109),
    .X(_06504_));
 sky130_fd_sc_hd__and4_1 _07204_ (.A(_06503_),
    .B(_06504_),
    .C(_05370_),
    .D(_05434_),
    .X(_06505_));
 sky130_fd_sc_hd__nor2_1 _07205_ (.A(_06502_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__xnor2_1 _07206_ (.A(_06499_),
    .B(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__nand3_1 _07207_ (.A(_06486_),
    .B(_06497_),
    .C(_06487_),
    .Y(_06508_));
 sky130_fd_sc_hd__a21bo_1 _07208_ (.A1(_06498_),
    .A2(_06507_),
    .B1_N(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__a21o_1 _07209_ (.A1(_06473_),
    .A2(_06474_),
    .B1(_06484_),
    .X(_06510_));
 sky130_fd_sc_hd__nand3_2 _07210_ (.A(_06485_),
    .B(_06509_),
    .C(_06510_),
    .Y(_06511_));
 sky130_fd_sc_hd__a21o_1 _07211_ (.A1(_06485_),
    .A2(_06510_),
    .B1(_06509_),
    .X(_06512_));
 sky130_fd_sc_hd__buf_4 _07212_ (.A(net66),
    .X(_06513_));
 sky130_fd_sc_hd__and4_1 _07213_ (.A(_02420_),
    .B(_06513_),
    .C(_05176_),
    .D(_05241_),
    .X(_06514_));
 sky130_fd_sc_hd__clkbuf_4 _07214_ (.A(net66),
    .X(_06515_));
 sky130_fd_sc_hd__buf_4 _07215_ (.A(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__buf_4 _07216_ (.A(_05176_),
    .X(_06517_));
 sky130_fd_sc_hd__buf_6 _07217_ (.A(net17),
    .X(_06518_));
 sky130_fd_sc_hd__clkbuf_4 _07218_ (.A(net107),
    .X(_06519_));
 sky130_fd_sc_hd__buf_4 _07219_ (.A(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__a22oi_1 _07220_ (.A1(_06516_),
    .A2(_06517_),
    .B1(_06518_),
    .B2(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__and4bb_1 _07221_ (.A_N(_06514_),
    .B_N(_06521_),
    .C(_02528_),
    .D(_05112_),
    .X(_06522_));
 sky130_fd_sc_hd__nor2_1 _07222_ (.A(_06514_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__o21ba_1 _07223_ (.A1(_06499_),
    .A2(_06502_),
    .B1_N(_06505_),
    .X(_06524_));
 sky130_fd_sc_hd__buf_4 _07224_ (.A(_05176_),
    .X(_06525_));
 sky130_fd_sc_hd__nand2_1 _07225_ (.A(_02528_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__and4_1 _07226_ (.A(_06519_),
    .B(_06515_),
    .C(net17),
    .D(net18),
    .X(_06527_));
 sky130_fd_sc_hd__a22o_1 _07227_ (.A1(_06515_),
    .A2(net17),
    .B1(_05305_),
    .B2(_06519_),
    .X(_06528_));
 sky130_fd_sc_hd__and2b_1 _07228_ (.A_N(_06527_),
    .B(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__xnor2_1 _07229_ (.A(_06526_),
    .B(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__xnor2_1 _07230_ (.A(_06524_),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__xnor2_1 _07231_ (.A(_06523_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand3_1 _07232_ (.A(_06511_),
    .B(_06512_),
    .C(_06532_),
    .Y(_06533_));
 sky130_fd_sc_hd__buf_6 _07233_ (.A(_02096_),
    .X(_06534_));
 sky130_fd_sc_hd__and4_1 _07234_ (.A(_06534_),
    .B(_06491_),
    .C(net130),
    .D(net129),
    .X(_06535_));
 sky130_fd_sc_hd__nand2_1 _07235_ (.A(_02248_),
    .B(_05638_),
    .Y(_06536_));
 sky130_fd_sc_hd__buf_4 _07236_ (.A(net130),
    .X(_06537_));
 sky130_fd_sc_hd__a22oi_4 _07237_ (.A1(_02205_),
    .A2(_06537_),
    .B1(_05756_),
    .B2(_02118_),
    .Y(_06538_));
 sky130_fd_sc_hd__or3_1 _07238_ (.A(_06535_),
    .B(_06536_),
    .C(_06538_),
    .X(_06539_));
 sky130_fd_sc_hd__o21bai_1 _07239_ (.A1(_06462_),
    .A2(_06464_),
    .B1_N(_06459_),
    .Y(_06540_));
 sky130_fd_sc_hd__o21ai_1 _07240_ (.A1(_06535_),
    .A2(_06538_),
    .B1(_06536_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand3_1 _07241_ (.A(_06539_),
    .B(_06540_),
    .C(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__a21o_1 _07242_ (.A1(_06539_),
    .A2(_06541_),
    .B1(_06540_),
    .X(_06543_));
 sky130_fd_sc_hd__buf_4 _07243_ (.A(net108),
    .X(_06544_));
 sky130_fd_sc_hd__buf_4 _07244_ (.A(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__buf_4 _07245_ (.A(_06489_),
    .X(_06546_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(_06545_),
    .B(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__buf_4 _07247_ (.A(net109),
    .X(_06548_));
 sky130_fd_sc_hd__and4_1 _07248_ (.A(_02291_),
    .B(_06548_),
    .C(_05498_),
    .D(_06461_),
    .X(_06549_));
 sky130_fd_sc_hd__a22o_1 _07249_ (.A1(_06548_),
    .A2(_05498_),
    .B1(_05563_),
    .B2(_02291_),
    .X(_06550_));
 sky130_fd_sc_hd__and2b_1 _07250_ (.A_N(_06549_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__xnor2_1 _07251_ (.A(_06547_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__nand3_1 _07252_ (.A(_06542_),
    .B(_06543_),
    .C(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__a21bo_1 _07253_ (.A1(_06474_),
    .A2(_06484_),
    .B1_N(_06473_),
    .X(_06554_));
 sky130_fd_sc_hd__a21o_1 _07254_ (.A1(_06542_),
    .A2(_06543_),
    .B1(_06552_),
    .X(_06555_));
 sky130_fd_sc_hd__nand3_2 _07255_ (.A(_06553_),
    .B(_06554_),
    .C(_06555_),
    .Y(_06556_));
 sky130_fd_sc_hd__a21o_1 _07256_ (.A1(_06553_),
    .A2(_06555_),
    .B1(_06554_),
    .X(_06557_));
 sky130_fd_sc_hd__a31o_1 _07257_ (.A1(_02550_),
    .A2(_05198_),
    .A3(_06528_),
    .B1(_06527_),
    .X(_06558_));
 sky130_fd_sc_hd__a31o_1 _07258_ (.A1(_02377_),
    .A2(_06477_),
    .A3(_06482_),
    .B1(_06481_),
    .X(_06559_));
 sky130_fd_sc_hd__buf_6 _07259_ (.A(net106),
    .X(_06560_));
 sky130_fd_sc_hd__clkbuf_8 _07260_ (.A(_06518_),
    .X(_06561_));
 sky130_fd_sc_hd__buf_4 _07261_ (.A(net18),
    .X(_06562_));
 sky130_fd_sc_hd__a22o_1 _07262_ (.A1(_06516_),
    .A2(_06562_),
    .B1(_06476_),
    .B2(_06520_),
    .X(_06563_));
 sky130_fd_sc_hd__buf_4 _07263_ (.A(net107),
    .X(_06564_));
 sky130_fd_sc_hd__clkbuf_4 _07264_ (.A(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__nand4_1 _07265_ (.A(_06565_),
    .B(_02485_),
    .C(_06562_),
    .D(_06476_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand4_1 _07266_ (.A(_06560_),
    .B(_06561_),
    .C(_06563_),
    .D(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__buf_4 _07267_ (.A(_05241_),
    .X(_06568_));
 sky130_fd_sc_hd__a22o_1 _07268_ (.A1(_06560_),
    .A2(_06568_),
    .B1(_06563_),
    .B2(_06566_),
    .X(_06569_));
 sky130_fd_sc_hd__and3_1 _07269_ (.A(_06559_),
    .B(_06567_),
    .C(_06569_),
    .X(_06570_));
 sky130_fd_sc_hd__a21o_1 _07270_ (.A1(_06567_),
    .A2(_06569_),
    .B1(_06559_),
    .X(_06571_));
 sky130_fd_sc_hd__and2b_1 _07271_ (.A_N(_06570_),
    .B(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__xor2_1 _07272_ (.A(_06558_),
    .B(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__a21oi_1 _07273_ (.A1(_06556_),
    .A2(_06557_),
    .B1(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__and3_1 _07274_ (.A(_06556_),
    .B(_06557_),
    .C(_06573_),
    .X(_06575_));
 sky130_fd_sc_hd__a211o_2 _07275_ (.A1(_06511_),
    .A2(_06533_),
    .B1(_06574_),
    .C1(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__o211ai_2 _07276_ (.A1(_06575_),
    .A2(_06574_),
    .B1(_06533_),
    .C1(_06511_),
    .Y(_06577_));
 sky130_fd_sc_hd__clkbuf_4 _07277_ (.A(net68),
    .X(_06578_));
 sky130_fd_sc_hd__clkbuf_4 _07278_ (.A(net38),
    .X(_06579_));
 sky130_fd_sc_hd__clkbuf_4 _07279_ (.A(net133),
    .X(_06580_));
 sky130_fd_sc_hd__clkbuf_4 _07280_ (.A(net13),
    .X(_06581_));
 sky130_fd_sc_hd__and4_1 _07281_ (.A(_06578_),
    .B(_06579_),
    .C(_06580_),
    .D(_06581_),
    .X(_06582_));
 sky130_fd_sc_hd__buf_4 _07282_ (.A(net38),
    .X(_06583_));
 sky130_fd_sc_hd__buf_4 _07283_ (.A(_06581_),
    .X(_06584_));
 sky130_fd_sc_hd__buf_4 _07284_ (.A(_02582_),
    .X(_06585_));
 sky130_fd_sc_hd__a22oi_1 _07285_ (.A1(_06583_),
    .A2(_04961_),
    .B1(_06584_),
    .B2(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__and4bb_1 _07286_ (.A_N(_06582_),
    .B_N(_06586_),
    .C(_02712_),
    .D(_04907_),
    .X(_06587_));
 sky130_fd_sc_hd__nor2_1 _07287_ (.A(_06582_),
    .B(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__and4_1 _07288_ (.A(_06578_),
    .B(_06579_),
    .C(_06581_),
    .D(_05101_),
    .X(_06589_));
 sky130_fd_sc_hd__a22oi_1 _07289_ (.A1(_06583_),
    .A2(_05025_),
    .B1(_05112_),
    .B2(_06585_),
    .Y(_06590_));
 sky130_fd_sc_hd__buf_4 _07290_ (.A(_06580_),
    .X(_06591_));
 sky130_fd_sc_hd__and4bb_1 _07291_ (.A_N(_06589_),
    .B_N(_06590_),
    .C(_02712_),
    .D(_06591_),
    .X(_06592_));
 sky130_fd_sc_hd__buf_4 _07292_ (.A(net122),
    .X(_06593_));
 sky130_fd_sc_hd__o2bb2a_1 _07293_ (.A1_N(_06593_),
    .A2_N(_04972_),
    .B1(_06589_),
    .B2(_06590_),
    .X(_06594_));
 sky130_fd_sc_hd__nor2_1 _07294_ (.A(_06592_),
    .B(_06594_),
    .Y(_06595_));
 sky130_fd_sc_hd__and2b_1 _07295_ (.A_N(_06588_),
    .B(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__xnor2_1 _07296_ (.A(_06588_),
    .B(_06595_),
    .Y(_06597_));
 sky130_fd_sc_hd__clkbuf_4 _07297_ (.A(net40),
    .X(_06598_));
 sky130_fd_sc_hd__clkbuf_4 _07298_ (.A(net41),
    .X(_06599_));
 sky130_fd_sc_hd__and4_1 _07299_ (.A(_06598_),
    .B(_06599_),
    .C(_04832_),
    .D(_04896_),
    .X(_06600_));
 sky130_fd_sc_hd__clkbuf_4 _07300_ (.A(net41),
    .X(_06601_));
 sky130_fd_sc_hd__buf_4 _07301_ (.A(net10),
    .X(_06602_));
 sky130_fd_sc_hd__clkbuf_8 _07302_ (.A(_06602_),
    .X(_06603_));
 sky130_fd_sc_hd__clkbuf_4 _07303_ (.A(net11),
    .X(_06604_));
 sky130_fd_sc_hd__buf_4 _07304_ (.A(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_4 _07305_ (.A(net40),
    .X(_06606_));
 sky130_fd_sc_hd__a22oi_1 _07306_ (.A1(_06601_),
    .A2(_06603_),
    .B1(_06605_),
    .B2(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__buf_4 _07307_ (.A(net121),
    .X(_06608_));
 sky130_fd_sc_hd__and4bb_1 _07308_ (.A_N(_06600_),
    .B_N(_06607_),
    .C(_06608_),
    .D(_04789_),
    .X(_06609_));
 sky130_fd_sc_hd__buf_6 _07309_ (.A(_06608_),
    .X(_06610_));
 sky130_fd_sc_hd__clkbuf_4 _07310_ (.A(net9),
    .X(_06611_));
 sky130_fd_sc_hd__buf_4 _07311_ (.A(_06611_),
    .X(_06612_));
 sky130_fd_sc_hd__buf_6 _07312_ (.A(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__o2bb2a_1 _07313_ (.A1_N(_06610_),
    .A2_N(_06613_),
    .B1(_06600_),
    .B2(_06607_),
    .X(_06614_));
 sky130_fd_sc_hd__nor2_1 _07314_ (.A(_06609_),
    .B(_06614_),
    .Y(_06615_));
 sky130_fd_sc_hd__and2_1 _07315_ (.A(_06597_),
    .B(_06615_),
    .X(_06616_));
 sky130_fd_sc_hd__or2b_1 _07316_ (.A(_06524_),
    .B_N(_06530_),
    .X(_06617_));
 sky130_fd_sc_hd__or2b_1 _07317_ (.A(_06523_),
    .B_N(_06531_),
    .X(_06618_));
 sky130_fd_sc_hd__nor2_1 _07318_ (.A(_06589_),
    .B(_06592_),
    .Y(_06619_));
 sky130_fd_sc_hd__buf_6 _07319_ (.A(net39),
    .X(_06620_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(_06620_),
    .B(_05047_),
    .Y(_06621_));
 sky130_fd_sc_hd__buf_4 _07321_ (.A(net38),
    .X(_06622_));
 sky130_fd_sc_hd__clkbuf_8 _07322_ (.A(net14),
    .X(_06623_));
 sky130_fd_sc_hd__and4_1 _07323_ (.A(_06585_),
    .B(_06622_),
    .C(_06623_),
    .D(_06517_),
    .X(_06624_));
 sky130_fd_sc_hd__a22o_1 _07324_ (.A1(_06583_),
    .A2(_06623_),
    .B1(_05187_),
    .B2(_06585_),
    .X(_06625_));
 sky130_fd_sc_hd__and2b_1 _07325_ (.A_N(_06624_),
    .B(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__xnor2_1 _07326_ (.A(_06621_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__xnor2_1 _07327_ (.A(_06619_),
    .B(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand2_4 _07328_ (.A(net121),
    .B(_04843_),
    .Y(_06629_));
 sky130_fd_sc_hd__buf_4 _07329_ (.A(_06599_),
    .X(_06630_));
 sky130_fd_sc_hd__buf_4 _07330_ (.A(_06598_),
    .X(_06631_));
 sky130_fd_sc_hd__a22oi_1 _07331_ (.A1(_06630_),
    .A2(_06605_),
    .B1(_06591_),
    .B2(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__and4_1 _07332_ (.A(_06598_),
    .B(_06599_),
    .C(_04896_),
    .D(_04961_),
    .X(_06633_));
 sky130_fd_sc_hd__nor2_1 _07333_ (.A(_06632_),
    .B(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__xnor2_2 _07334_ (.A(_06629_),
    .B(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__xnor2_1 _07335_ (.A(_06628_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__a21o_2 _07336_ (.A1(_06617_),
    .A2(_06618_),
    .B1(_06636_),
    .X(_06637_));
 sky130_fd_sc_hd__nand3_1 _07337_ (.A(_06617_),
    .B(_06618_),
    .C(_06636_),
    .Y(_06638_));
 sky130_fd_sc_hd__o211ai_4 _07338_ (.A1(_06596_),
    .A2(_06616_),
    .B1(_06637_),
    .C1(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__a211o_1 _07339_ (.A1(_06637_),
    .A2(_06638_),
    .B1(_06596_),
    .C1(_06616_),
    .X(_06640_));
 sky130_fd_sc_hd__nand4_4 _07340_ (.A(_06576_),
    .B(_06577_),
    .C(_06639_),
    .D(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nand3_1 _07341_ (.A(_06556_),
    .B(_06557_),
    .C(_06573_),
    .Y(_06642_));
 sky130_fd_sc_hd__and4_1 _07342_ (.A(_02107_),
    .B(_06495_),
    .C(net129),
    .D(net128),
    .X(_06643_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_02248_),
    .B(net130),
    .Y(_06644_));
 sky130_fd_sc_hd__a22oi_2 _07344_ (.A1(_02205_),
    .A2(net129),
    .B1(net128),
    .B2(_06534_),
    .Y(_06645_));
 sky130_fd_sc_hd__or3_1 _07345_ (.A(_06643_),
    .B(_06644_),
    .C(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__o21bai_1 _07346_ (.A1(_06536_),
    .A2(_06538_),
    .B1_N(_06535_),
    .Y(_06647_));
 sky130_fd_sc_hd__o21ai_1 _07347_ (.A1(_06643_),
    .A2(_06645_),
    .B1(_06644_),
    .Y(_06648_));
 sky130_fd_sc_hd__nand3_1 _07348_ (.A(_06646_),
    .B(_06647_),
    .C(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__a21o_1 _07349_ (.A1(_06646_),
    .A2(_06648_),
    .B1(_06647_),
    .X(_06650_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(_06544_),
    .B(_05498_),
    .Y(_06651_));
 sky130_fd_sc_hd__and4_1 _07351_ (.A(_06479_),
    .B(_06480_),
    .C(_06461_),
    .D(_05627_),
    .X(_06652_));
 sky130_fd_sc_hd__a22oi_1 _07352_ (.A1(_06500_),
    .A2(_05563_),
    .B1(_05638_),
    .B2(_06501_),
    .Y(_06653_));
 sky130_fd_sc_hd__nor2_1 _07353_ (.A(_06652_),
    .B(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__xnor2_1 _07354_ (.A(_06651_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__nand3_1 _07355_ (.A(_06649_),
    .B(_06650_),
    .C(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__a21bo_1 _07356_ (.A1(_06543_),
    .A2(_06552_),
    .B1_N(_06542_),
    .X(_06657_));
 sky130_fd_sc_hd__a21o_1 _07357_ (.A1(_06649_),
    .A2(_06650_),
    .B1(_06655_),
    .X(_06658_));
 sky130_fd_sc_hd__nand3_2 _07358_ (.A(_06656_),
    .B(_06657_),
    .C(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__a21o_1 _07359_ (.A1(_06656_),
    .A2(_06658_),
    .B1(_06657_),
    .X(_06660_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(_06566_),
    .B(_06567_),
    .Y(_06661_));
 sky130_fd_sc_hd__a31o_1 _07361_ (.A1(_02377_),
    .A2(_06546_),
    .A3(_06550_),
    .B1(_06549_),
    .X(_06662_));
 sky130_fd_sc_hd__buf_4 _07362_ (.A(net106),
    .X(_06663_));
 sky130_fd_sc_hd__nand2_1 _07363_ (.A(_06663_),
    .B(_05316_),
    .Y(_06664_));
 sky130_fd_sc_hd__a22o_1 _07364_ (.A1(_06516_),
    .A2(_05370_),
    .B1(_06489_),
    .B2(_06520_),
    .X(_06665_));
 sky130_fd_sc_hd__buf_4 _07365_ (.A(_05434_),
    .X(_06666_));
 sky130_fd_sc_hd__nand4_1 _07366_ (.A(_06565_),
    .B(_02485_),
    .C(_06476_),
    .D(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand3b_1 _07367_ (.A_N(_06664_),
    .B(_06665_),
    .C(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__a21bo_1 _07368_ (.A1(_06665_),
    .A2(_06667_),
    .B1_N(_06664_),
    .X(_06669_));
 sky130_fd_sc_hd__and3_1 _07369_ (.A(_06662_),
    .B(_06668_),
    .C(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a21o_1 _07370_ (.A1(_06668_),
    .A2(_06669_),
    .B1(_06662_),
    .X(_06671_));
 sky130_fd_sc_hd__and2b_1 _07371_ (.A_N(_06670_),
    .B(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__xor2_1 _07372_ (.A(_06661_),
    .B(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__a21oi_2 _07373_ (.A1(_06659_),
    .A2(_06660_),
    .B1(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__and3_1 _07374_ (.A(_06659_),
    .B(_06660_),
    .C(_06673_),
    .X(_06675_));
 sky130_fd_sc_hd__a211oi_4 _07375_ (.A1(_06556_),
    .A2(_06642_),
    .B1(_06674_),
    .C1(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__o211a_1 _07376_ (.A1(_06675_),
    .A2(_06674_),
    .B1(_06642_),
    .C1(_06556_),
    .X(_06677_));
 sky130_fd_sc_hd__and2b_1 _07377_ (.A_N(_06619_),
    .B(_06627_),
    .X(_06678_));
 sky130_fd_sc_hd__and2_1 _07378_ (.A(_06628_),
    .B(_06635_),
    .X(_06679_));
 sky130_fd_sc_hd__buf_4 _07379_ (.A(net39),
    .X(_06680_));
 sky130_fd_sc_hd__and2_1 _07380_ (.A(_06680_),
    .B(_05112_),
    .X(_06681_));
 sky130_fd_sc_hd__buf_4 _07381_ (.A(_06579_),
    .X(_06682_));
 sky130_fd_sc_hd__buf_4 _07382_ (.A(_06578_),
    .X(_00000_));
 sky130_fd_sc_hd__a22o_1 _07383_ (.A1(_06682_),
    .A2(_06525_),
    .B1(_06568_),
    .B2(_00000_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_4 _07384_ (.A(_06517_),
    .X(_00002_));
 sky130_fd_sc_hd__nand4_1 _07385_ (.A(_00000_),
    .B(_06682_),
    .C(_00002_),
    .D(_06568_),
    .Y(_00003_));
 sky130_fd_sc_hd__nand3_1 _07386_ (.A(_06681_),
    .B(_00001_),
    .C(_00003_),
    .Y(_00004_));
 sky130_fd_sc_hd__a21o_1 _07387_ (.A1(_00001_),
    .A2(_00003_),
    .B1(_06681_),
    .X(_00005_));
 sky130_fd_sc_hd__a31o_1 _07388_ (.A1(_02723_),
    .A2(_05047_),
    .A3(_06625_),
    .B1(_06624_),
    .X(_00006_));
 sky130_fd_sc_hd__nand3_1 _07389_ (.A(_00004_),
    .B(_00005_),
    .C(_00006_),
    .Y(_00007_));
 sky130_fd_sc_hd__a21o_1 _07390_ (.A1(_00004_),
    .A2(_00005_),
    .B1(_00006_),
    .X(_00008_));
 sky130_fd_sc_hd__nand2_1 _07391_ (.A(_02851_),
    .B(_04918_),
    .Y(_00009_));
 sky130_fd_sc_hd__and3_1 _07392_ (.A(_06606_),
    .B(_06601_),
    .C(_06584_),
    .X(_00010_));
 sky130_fd_sc_hd__buf_6 _07393_ (.A(_06599_),
    .X(_00011_));
 sky130_fd_sc_hd__buf_6 _07394_ (.A(_06598_),
    .X(_00012_));
 sky130_fd_sc_hd__a22o_1 _07395_ (.A1(_00011_),
    .A2(_06591_),
    .B1(_05036_),
    .B2(_00012_),
    .X(_00013_));
 sky130_fd_sc_hd__a21bo_1 _07396_ (.A1(_04983_),
    .A2(_00010_),
    .B1_N(_00013_),
    .X(_00014_));
 sky130_fd_sc_hd__xor2_1 _07397_ (.A(_00009_),
    .B(_00014_),
    .X(_00015_));
 sky130_fd_sc_hd__nand3_1 _07398_ (.A(_00007_),
    .B(_00008_),
    .C(_00015_),
    .Y(_00016_));
 sky130_fd_sc_hd__a21o_1 _07399_ (.A1(_00007_),
    .A2(_00008_),
    .B1(_00015_),
    .X(_00017_));
 sky130_fd_sc_hd__a21o_1 _07400_ (.A1(_06558_),
    .A2(_06571_),
    .B1(_06570_),
    .X(_00018_));
 sky130_fd_sc_hd__a21o_1 _07401_ (.A1(_00016_),
    .A2(_00017_),
    .B1(_00018_),
    .X(_00019_));
 sky130_fd_sc_hd__nand3_1 _07402_ (.A(_00018_),
    .B(_00016_),
    .C(_00017_),
    .Y(_00020_));
 sky130_fd_sc_hd__o211ai_2 _07403_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_00019_),
    .C1(_00020_),
    .Y(_00021_));
 sky130_fd_sc_hd__a211o_1 _07404_ (.A1(_00020_),
    .A2(_00019_),
    .B1(_06679_),
    .C1(_06678_),
    .X(_00022_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(_00021_),
    .B(_00022_),
    .Y(_00023_));
 sky130_fd_sc_hd__o21a_1 _07406_ (.A1(_06676_),
    .A2(_06677_),
    .B1(_00023_),
    .X(_00024_));
 sky130_fd_sc_hd__nor3_4 _07407_ (.A(_06676_),
    .B(_06677_),
    .C(_00023_),
    .Y(_00025_));
 sky130_fd_sc_hd__a211o_1 _07408_ (.A1(_06576_),
    .A2(_06641_),
    .B1(_00024_),
    .C1(_00025_),
    .X(_00026_));
 sky130_fd_sc_hd__o211ai_2 _07409_ (.A1(_00025_),
    .A2(_00024_),
    .B1(_06641_),
    .C1(_06576_),
    .Y(_00027_));
 sky130_fd_sc_hd__clkbuf_4 _07410_ (.A(net120),
    .X(_00028_));
 sky130_fd_sc_hd__buf_4 _07411_ (.A(net44),
    .X(_00029_));
 sky130_fd_sc_hd__clkbuf_4 _07412_ (.A(net7),
    .X(_00030_));
 sky130_fd_sc_hd__and4_1 _07413_ (.A(_00028_),
    .B(_00029_),
    .C(_00030_),
    .D(_04703_),
    .X(_00031_));
 sky130_fd_sc_hd__clkbuf_4 _07414_ (.A(net8),
    .X(_00032_));
 sky130_fd_sc_hd__buf_4 _07415_ (.A(_00032_),
    .X(_00033_));
 sky130_fd_sc_hd__a22oi_1 _07416_ (.A1(_02948_),
    .A2(_04638_),
    .B1(_00033_),
    .B2(_02894_),
    .Y(_00034_));
 sky130_fd_sc_hd__buf_4 _07417_ (.A(net6),
    .X(_00035_));
 sky130_fd_sc_hd__buf_4 _07418_ (.A(_00035_),
    .X(_00036_));
 sky130_fd_sc_hd__and4bb_1 _07419_ (.A_N(_00031_),
    .B_N(_00034_),
    .C(net119),
    .D(_00036_),
    .X(_00037_));
 sky130_fd_sc_hd__and4_1 _07420_ (.A(net40),
    .B(net41),
    .C(_06611_),
    .D(_06602_),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _07421_ (.A1(_06599_),
    .A2(_06611_),
    .B1(_04832_),
    .B2(_06598_),
    .X(_00039_));
 sky130_fd_sc_hd__buf_6 _07422_ (.A(_04703_),
    .X(_00040_));
 sky130_fd_sc_hd__and4b_1 _07423_ (.A_N(_00038_),
    .B(_00039_),
    .C(net121),
    .D(_00040_),
    .X(_00041_));
 sky130_fd_sc_hd__nor2_1 _07424_ (.A(_00038_),
    .B(_00041_),
    .Y(_00042_));
 sky130_fd_sc_hd__o2bb2a_1 _07425_ (.A1_N(_03002_),
    .A2_N(_00036_),
    .B1(_00031_),
    .B2(_00034_),
    .X(_00043_));
 sky130_fd_sc_hd__or3_1 _07426_ (.A(_00037_),
    .B(_00042_),
    .C(_00043_),
    .X(_00044_));
 sky130_fd_sc_hd__and4_1 _07427_ (.A(_00028_),
    .B(_00029_),
    .C(_00035_),
    .D(_04638_),
    .X(_00045_));
 sky130_fd_sc_hd__buf_4 _07428_ (.A(net44),
    .X(_00046_));
 sky130_fd_sc_hd__buf_4 _07429_ (.A(_04574_),
    .X(_00047_));
 sky130_fd_sc_hd__buf_4 _07430_ (.A(_00030_),
    .X(_00048_));
 sky130_fd_sc_hd__buf_6 _07431_ (.A(net43),
    .X(_00049_));
 sky130_fd_sc_hd__a22oi_2 _07432_ (.A1(_00046_),
    .A2(_00047_),
    .B1(_00048_),
    .B2(_00049_),
    .Y(_00050_));
 sky130_fd_sc_hd__and4bb_1 _07433_ (.A_N(_00045_),
    .B_N(_00050_),
    .C(_03002_),
    .D(_04520_),
    .X(_00051_));
 sky130_fd_sc_hd__or2_1 _07434_ (.A(_00045_),
    .B(_00051_),
    .X(_00052_));
 sky130_fd_sc_hd__nor2_1 _07435_ (.A(_00037_),
    .B(_00043_),
    .Y(_00053_));
 sky130_fd_sc_hd__xnor2_1 _07436_ (.A(_00042_),
    .B(_00053_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand2_1 _07437_ (.A(_00052_),
    .B(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__or2_1 _07438_ (.A(_00031_),
    .B(_00037_),
    .X(_00056_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_06600_),
    .B(_06609_),
    .Y(_00057_));
 sky130_fd_sc_hd__buf_6 _07440_ (.A(net119),
    .X(_00058_));
 sky130_fd_sc_hd__buf_6 _07441_ (.A(_00048_),
    .X(_00059_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(_00058_),
    .B(_00059_),
    .Y(_00060_));
 sky130_fd_sc_hd__and4_1 _07443_ (.A(_02894_),
    .B(_02948_),
    .C(_04703_),
    .D(_04778_),
    .X(_00061_));
 sky130_fd_sc_hd__buf_6 _07444_ (.A(_00029_),
    .X(_00062_));
 sky130_fd_sc_hd__buf_4 _07445_ (.A(_00028_),
    .X(_00063_));
 sky130_fd_sc_hd__a22oi_1 _07446_ (.A1(_00062_),
    .A2(_00040_),
    .B1(_06612_),
    .B2(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__nor2_1 _07447_ (.A(_00061_),
    .B(_00064_),
    .Y(_00065_));
 sky130_fd_sc_hd__xnor2_1 _07448_ (.A(_00060_),
    .B(_00065_),
    .Y(_00066_));
 sky130_fd_sc_hd__xnor2_1 _07449_ (.A(_00057_),
    .B(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__xnor2_1 _07450_ (.A(_00056_),
    .B(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__a21o_1 _07451_ (.A1(_00044_),
    .A2(_00055_),
    .B1(_00068_),
    .X(_00069_));
 sky130_fd_sc_hd__a21oi_1 _07452_ (.A1(_00044_),
    .A2(_00055_),
    .B1(_00068_),
    .Y(_00070_));
 sky130_fd_sc_hd__and3_1 _07453_ (.A(_00044_),
    .B(_00055_),
    .C(_00068_),
    .X(_00071_));
 sky130_fd_sc_hd__buf_4 _07454_ (.A(net34),
    .X(_00072_));
 sky130_fd_sc_hd__and4_1 _07455_ (.A(net50),
    .B(net51),
    .C(_04294_),
    .D(_00072_),
    .X(_00073_));
 sky130_fd_sc_hd__clkbuf_4 _07456_ (.A(net123),
    .X(_00074_));
 sky130_fd_sc_hd__a22oi_1 _07457_ (.A1(_03271_),
    .A2(_00074_),
    .B1(_04358_),
    .B2(_03217_),
    .Y(_00075_));
 sky130_fd_sc_hd__and4bb_1 _07458_ (.A_N(_00073_),
    .B_N(_00075_),
    .C(net114),
    .D(_04240_),
    .X(_00076_));
 sky130_fd_sc_hd__buf_4 _07459_ (.A(net114),
    .X(_00077_));
 sky130_fd_sc_hd__o2bb2a_1 _07460_ (.A1_N(_00077_),
    .A2_N(_04251_),
    .B1(_00073_),
    .B2(_00075_),
    .X(_00078_));
 sky130_fd_sc_hd__nor2_1 _07461_ (.A(_00076_),
    .B(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__and4_1 _07462_ (.A(net118),
    .B(net117),
    .C(_04434_),
    .D(_04509_),
    .X(_00080_));
 sky130_fd_sc_hd__clkbuf_4 _07463_ (.A(net117),
    .X(_00081_));
 sky130_fd_sc_hd__buf_2 _07464_ (.A(net35),
    .X(_00082_));
 sky130_fd_sc_hd__buf_4 _07465_ (.A(_00082_),
    .X(_00083_));
 sky130_fd_sc_hd__buf_2 _07466_ (.A(net36),
    .X(_00084_));
 sky130_fd_sc_hd__buf_4 _07467_ (.A(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__buf_4 _07468_ (.A(net118),
    .X(_00086_));
 sky130_fd_sc_hd__a22oi_1 _07469_ (.A1(_00081_),
    .A2(_00083_),
    .B1(_00085_),
    .B2(_00086_),
    .Y(_00087_));
 sky130_fd_sc_hd__buf_6 _07470_ (.A(net49),
    .X(_00088_));
 sky130_fd_sc_hd__buf_4 _07471_ (.A(net34),
    .X(_00089_));
 sky130_fd_sc_hd__buf_4 _07472_ (.A(_00089_),
    .X(_00090_));
 sky130_fd_sc_hd__and4bb_1 _07473_ (.A_N(_00080_),
    .B_N(_00087_),
    .C(_00088_),
    .D(_00090_),
    .X(_00091_));
 sky130_fd_sc_hd__nor2_1 _07474_ (.A(_00080_),
    .B(_00091_),
    .Y(_00092_));
 sky130_fd_sc_hd__buf_6 _07475_ (.A(_04434_),
    .X(_00093_));
 sky130_fd_sc_hd__nand2_1 _07476_ (.A(_03163_),
    .B(_00093_),
    .Y(_00094_));
 sky130_fd_sc_hd__buf_2 _07477_ (.A(net118),
    .X(_00095_));
 sky130_fd_sc_hd__clkbuf_4 _07478_ (.A(net117),
    .X(_00096_));
 sky130_fd_sc_hd__and4_1 _07479_ (.A(_00095_),
    .B(_00096_),
    .C(_04509_),
    .D(_00035_),
    .X(_00097_));
 sky130_fd_sc_hd__buf_4 _07480_ (.A(_00084_),
    .X(_00098_));
 sky130_fd_sc_hd__a22oi_1 _07481_ (.A1(_03099_),
    .A2(_00098_),
    .B1(_00047_),
    .B2(_03056_),
    .Y(_00099_));
 sky130_fd_sc_hd__nor2_1 _07482_ (.A(_00097_),
    .B(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__xnor2_1 _07483_ (.A(_00094_),
    .B(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__xnor2_1 _07484_ (.A(_00092_),
    .B(_00101_),
    .Y(_00102_));
 sky130_fd_sc_hd__and2_1 _07485_ (.A(_00079_),
    .B(_00102_),
    .X(_00103_));
 sky130_fd_sc_hd__nor2_1 _07486_ (.A(_00079_),
    .B(_00102_),
    .Y(_00104_));
 sky130_fd_sc_hd__or2_2 _07487_ (.A(_00103_),
    .B(_00104_),
    .X(_00105_));
 sky130_fd_sc_hd__or3_1 _07488_ (.A(_00070_),
    .B(_00071_),
    .C(_00105_),
    .X(_00106_));
 sky130_fd_sc_hd__or2b_1 _07489_ (.A(_00057_),
    .B_N(_00066_),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(_00056_),
    .B(_00067_),
    .Y(_00108_));
 sky130_fd_sc_hd__and4_1 _07491_ (.A(net120),
    .B(net44),
    .C(_06611_),
    .D(_06602_),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(net119),
    .B(_00033_),
    .Y(_00110_));
 sky130_fd_sc_hd__a22oi_1 _07493_ (.A1(_02948_),
    .A2(_04778_),
    .B1(_06603_),
    .B2(_02894_),
    .Y(_00111_));
 sky130_fd_sc_hd__or3_1 _07494_ (.A(_00109_),
    .B(_00110_),
    .C(_00111_),
    .X(_00112_));
 sky130_fd_sc_hd__o21bai_1 _07495_ (.A1(_06629_),
    .A2(_06632_),
    .B1_N(_06633_),
    .Y(_00113_));
 sky130_fd_sc_hd__o21ai_1 _07496_ (.A1(_00109_),
    .A2(_00111_),
    .B1(_00110_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand3_1 _07497_ (.A(_00112_),
    .B(_00113_),
    .C(_00114_),
    .Y(_00115_));
 sky130_fd_sc_hd__a31o_1 _07498_ (.A1(_03013_),
    .A2(_04660_),
    .A3(_00065_),
    .B1(_00061_),
    .X(_00116_));
 sky130_fd_sc_hd__a21o_1 _07499_ (.A1(_00112_),
    .A2(_00114_),
    .B1(_00113_),
    .X(_00117_));
 sky130_fd_sc_hd__and3_1 _07500_ (.A(_00115_),
    .B(_00116_),
    .C(_00117_),
    .X(_00118_));
 sky130_fd_sc_hd__a21oi_1 _07501_ (.A1(_00115_),
    .A2(_00117_),
    .B1(_00116_),
    .Y(_00119_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(_00118_),
    .B(_00119_),
    .X(_00120_));
 sky130_fd_sc_hd__a21oi_4 _07503_ (.A1(_00107_),
    .A2(_00108_),
    .B1(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__and3_1 _07504_ (.A(_00107_),
    .B(_00108_),
    .C(_00120_),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_2 _07505_ (.A(_00077_),
    .B(_04316_),
    .Y(_00123_));
 sky130_fd_sc_hd__buf_4 _07506_ (.A(net50),
    .X(_00124_));
 sky130_fd_sc_hd__buf_4 _07507_ (.A(net51),
    .X(_00125_));
 sky130_fd_sc_hd__and3_1 _07508_ (.A(_00124_),
    .B(_00125_),
    .C(_04445_),
    .X(_00126_));
 sky130_fd_sc_hd__a22o_1 _07509_ (.A1(_00125_),
    .A2(_00090_),
    .B1(_04445_),
    .B2(_00124_),
    .X(_00127_));
 sky130_fd_sc_hd__a21bo_1 _07510_ (.A1(_04369_),
    .A2(_00126_),
    .B1_N(_00127_),
    .X(_00128_));
 sky130_fd_sc_hd__xor2_4 _07511_ (.A(_00123_),
    .B(_00128_),
    .X(_00129_));
 sky130_fd_sc_hd__and4_1 _07512_ (.A(_00086_),
    .B(_00081_),
    .C(_00047_),
    .D(_04638_),
    .X(_00130_));
 sky130_fd_sc_hd__nand2_1 _07513_ (.A(_00088_),
    .B(_04520_),
    .Y(_00131_));
 sky130_fd_sc_hd__buf_4 _07514_ (.A(net117),
    .X(_00132_));
 sky130_fd_sc_hd__buf_4 _07515_ (.A(net118),
    .X(_00133_));
 sky130_fd_sc_hd__a22oi_2 _07516_ (.A1(_00132_),
    .A2(_00047_),
    .B1(_00048_),
    .B2(_00133_),
    .Y(_00134_));
 sky130_fd_sc_hd__or3_1 _07517_ (.A(_00130_),
    .B(_00131_),
    .C(_00134_),
    .X(_00135_));
 sky130_fd_sc_hd__o21ai_1 _07518_ (.A1(_00130_),
    .A2(_00134_),
    .B1(_00131_),
    .Y(_00136_));
 sky130_fd_sc_hd__o21bai_1 _07519_ (.A1(_00094_),
    .A2(_00099_),
    .B1_N(_00097_),
    .Y(_00137_));
 sky130_fd_sc_hd__and3_1 _07520_ (.A(_00135_),
    .B(_00136_),
    .C(_00137_),
    .X(_00138_));
 sky130_fd_sc_hd__a21o_1 _07521_ (.A1(_00135_),
    .A2(_00136_),
    .B1(_00137_),
    .X(_00139_));
 sky130_fd_sc_hd__and2b_1 _07522_ (.A_N(_00138_),
    .B(_00139_),
    .X(_00140_));
 sky130_fd_sc_hd__xnor2_4 _07523_ (.A(_00129_),
    .B(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__o21a_1 _07524_ (.A1(_00121_),
    .A2(_00122_),
    .B1(_00141_),
    .X(_00142_));
 sky130_fd_sc_hd__nor3_4 _07525_ (.A(_00121_),
    .B(_00122_),
    .C(_00141_),
    .Y(_00143_));
 sky130_fd_sc_hd__a211oi_4 _07526_ (.A1(_06637_),
    .A2(_06639_),
    .B1(_00142_),
    .C1(_00143_),
    .Y(_00144_));
 sky130_fd_sc_hd__o211a_1 _07527_ (.A1(_00143_),
    .A2(_00142_),
    .B1(_06639_),
    .C1(_06637_),
    .X(_00145_));
 sky130_fd_sc_hd__a211o_1 _07528_ (.A1(_00069_),
    .A2(_00106_),
    .B1(_00144_),
    .C1(_00145_),
    .X(_00146_));
 sky130_fd_sc_hd__o211ai_2 _07529_ (.A1(_00144_),
    .A2(_00145_),
    .B1(_00069_),
    .C1(_00106_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand4_1 _07530_ (.A(_00026_),
    .B(_00027_),
    .C(_00146_),
    .D(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand3_1 _07531_ (.A(_06659_),
    .B(_06660_),
    .C(_06673_),
    .Y(_00149_));
 sky130_fd_sc_hd__buf_4 _07532_ (.A(net116),
    .X(_00150_));
 sky130_fd_sc_hd__and4_1 _07533_ (.A(_06494_),
    .B(_00150_),
    .C(net128),
    .D(net28),
    .X(_00151_));
 sky130_fd_sc_hd__nand2_1 _07534_ (.A(_06488_),
    .B(net129),
    .Y(_00152_));
 sky130_fd_sc_hd__clkbuf_4 _07535_ (.A(net28),
    .X(_00153_));
 sky130_fd_sc_hd__a22oi_2 _07536_ (.A1(_06491_),
    .A2(net128),
    .B1(_00153_),
    .B2(_06492_),
    .Y(_00154_));
 sky130_fd_sc_hd__or3_1 _07537_ (.A(_00151_),
    .B(_00152_),
    .C(_00154_),
    .X(_00155_));
 sky130_fd_sc_hd__o21bai_1 _07538_ (.A1(_06644_),
    .A2(_06645_),
    .B1_N(_06643_),
    .Y(_00156_));
 sky130_fd_sc_hd__o21ai_1 _07539_ (.A1(_00151_),
    .A2(_00154_),
    .B1(_00152_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand3_1 _07540_ (.A(_00155_),
    .B(_00156_),
    .C(_00157_),
    .Y(_00158_));
 sky130_fd_sc_hd__a21o_1 _07541_ (.A1(_00155_),
    .A2(_00157_),
    .B1(_00156_),
    .X(_00159_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(_06475_),
    .B(_05574_),
    .Y(_00160_));
 sky130_fd_sc_hd__and4_1 _07543_ (.A(_02291_),
    .B(_06548_),
    .C(_05627_),
    .D(net130),
    .X(_00161_));
 sky130_fd_sc_hd__buf_4 _07544_ (.A(_06480_),
    .X(_00162_));
 sky130_fd_sc_hd__clkbuf_4 _07545_ (.A(net130),
    .X(_00163_));
 sky130_fd_sc_hd__buf_4 _07546_ (.A(_06479_),
    .X(_00164_));
 sky130_fd_sc_hd__a22oi_1 _07547_ (.A1(_00162_),
    .A2(_05638_),
    .B1(_00163_),
    .B2(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__nor2_1 _07548_ (.A(_00161_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__xnor2_1 _07549_ (.A(_00160_),
    .B(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand3_1 _07550_ (.A(_00158_),
    .B(_00159_),
    .C(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__a21bo_1 _07551_ (.A1(_06650_),
    .A2(_06655_),
    .B1_N(_06649_),
    .X(_00169_));
 sky130_fd_sc_hd__a21o_1 _07552_ (.A1(_00158_),
    .A2(_00159_),
    .B1(_00167_),
    .X(_00170_));
 sky130_fd_sc_hd__nand3_1 _07553_ (.A(_00168_),
    .B(_00169_),
    .C(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__a21o_1 _07554_ (.A1(_00168_),
    .A2(_00170_),
    .B1(_00169_),
    .X(_00172_));
 sky130_fd_sc_hd__nand2_1 _07555_ (.A(_06667_),
    .B(_06668_),
    .Y(_00173_));
 sky130_fd_sc_hd__o21bai_1 _07556_ (.A1(_06651_),
    .A2(_06653_),
    .B1_N(_06652_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(net106),
    .B(_06476_),
    .Y(_00175_));
 sky130_fd_sc_hd__a22o_1 _07558_ (.A1(_06513_),
    .A2(_05434_),
    .B1(_06466_),
    .B2(_02420_),
    .X(_00176_));
 sky130_fd_sc_hd__nand4_1 _07559_ (.A(_02420_),
    .B(_06513_),
    .C(_05434_),
    .D(_06466_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand3b_1 _07560_ (.A_N(_00175_),
    .B(_00176_),
    .C(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__a21bo_1 _07561_ (.A1(_00176_),
    .A2(_00177_),
    .B1_N(_00175_),
    .X(_00179_));
 sky130_fd_sc_hd__and3_1 _07562_ (.A(_00174_),
    .B(_00178_),
    .C(_00179_),
    .X(_00180_));
 sky130_fd_sc_hd__a21o_1 _07563_ (.A1(_00178_),
    .A2(_00179_),
    .B1(_00174_),
    .X(_00181_));
 sky130_fd_sc_hd__and2b_1 _07564_ (.A_N(_00180_),
    .B(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__xor2_1 _07565_ (.A(_00173_),
    .B(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__a21oi_2 _07566_ (.A1(_00171_),
    .A2(_00172_),
    .B1(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__and3_2 _07567_ (.A(_00171_),
    .B(_00172_),
    .C(_00183_),
    .X(_00185_));
 sky130_fd_sc_hd__a211oi_4 _07568_ (.A1(_06659_),
    .A2(_00149_),
    .B1(_00184_),
    .C1(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__o211a_1 _07569_ (.A1(_00185_),
    .A2(_00184_),
    .B1(_00149_),
    .C1(_06659_),
    .X(_00187_));
 sky130_fd_sc_hd__a21o_1 _07570_ (.A1(_06661_),
    .A2(_06671_),
    .B1(_06670_),
    .X(_00188_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(_06680_),
    .B(_06525_),
    .Y(_00189_));
 sky130_fd_sc_hd__a22oi_2 _07572_ (.A1(_02658_),
    .A2(_05252_),
    .B1(_05316_),
    .B2(_02593_),
    .Y(_00190_));
 sky130_fd_sc_hd__and4_1 _07573_ (.A(_06585_),
    .B(_06583_),
    .C(_06518_),
    .D(_06562_),
    .X(_00191_));
 sky130_fd_sc_hd__or3_1 _07574_ (.A(_00189_),
    .B(_00190_),
    .C(_00191_),
    .X(_00192_));
 sky130_fd_sc_hd__o21ai_1 _07575_ (.A1(_00190_),
    .A2(_00191_),
    .B1(_00189_),
    .Y(_00193_));
 sky130_fd_sc_hd__a21bo_1 _07576_ (.A1(_06681_),
    .A2(_00001_),
    .B1_N(_00003_),
    .X(_00194_));
 sky130_fd_sc_hd__nand3_1 _07577_ (.A(_00192_),
    .B(_00193_),
    .C(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__a21o_1 _07578_ (.A1(_00192_),
    .A2(_00193_),
    .B1(_00194_),
    .X(_00196_));
 sky130_fd_sc_hd__buf_4 _07579_ (.A(_04961_),
    .X(_00197_));
 sky130_fd_sc_hd__nand2_1 _07580_ (.A(_06610_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__a22o_1 _07581_ (.A1(_06601_),
    .A2(_06584_),
    .B1(_05112_),
    .B2(_06606_),
    .X(_00199_));
 sky130_fd_sc_hd__a21bo_1 _07582_ (.A1(_05123_),
    .A2(_00010_),
    .B1_N(_00199_),
    .X(_00200_));
 sky130_fd_sc_hd__xor2_1 _07583_ (.A(_00198_),
    .B(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__nand3_1 _07584_ (.A(_00195_),
    .B(_00196_),
    .C(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__a21o_1 _07585_ (.A1(_00195_),
    .A2(_00196_),
    .B1(_00201_),
    .X(_00203_));
 sky130_fd_sc_hd__nand3_1 _07586_ (.A(_00188_),
    .B(_00202_),
    .C(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _07587_ (.A(_00007_),
    .B(_00016_),
    .Y(_00205_));
 sky130_fd_sc_hd__a21o_1 _07588_ (.A1(_00202_),
    .A2(_00203_),
    .B1(_00188_),
    .X(_00206_));
 sky130_fd_sc_hd__nand3_1 _07589_ (.A(_00204_),
    .B(_00205_),
    .C(_00206_),
    .Y(_00207_));
 sky130_fd_sc_hd__a21o_1 _07590_ (.A1(_00204_),
    .A2(_00206_),
    .B1(_00205_),
    .X(_00208_));
 sky130_fd_sc_hd__nand2_1 _07591_ (.A(_00207_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__o21ai_2 _07592_ (.A1(_00186_),
    .A2(_00187_),
    .B1(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__or3_1 _07593_ (.A(_00186_),
    .B(_00187_),
    .C(_00209_),
    .X(_00211_));
 sky130_fd_sc_hd__o211ai_4 _07594_ (.A1(_06676_),
    .A2(_00025_),
    .B1(_00210_),
    .C1(_00211_),
    .Y(_00212_));
 sky130_fd_sc_hd__a211o_1 _07595_ (.A1(_00211_),
    .A2(_00210_),
    .B1(_00025_),
    .C1(_06676_),
    .X(_00213_));
 sky130_fd_sc_hd__or2b_1 _07596_ (.A(_00109_),
    .B_N(_00112_),
    .X(_00214_));
 sky130_fd_sc_hd__a32o_1 _07597_ (.A1(_06610_),
    .A2(_04918_),
    .A3(_00013_),
    .B1(_00010_),
    .B2(_00197_),
    .X(_00215_));
 sky130_fd_sc_hd__buf_4 _07598_ (.A(_00029_),
    .X(_00216_));
 sky130_fd_sc_hd__buf_4 _07599_ (.A(_00028_),
    .X(_00217_));
 sky130_fd_sc_hd__a22o_1 _07600_ (.A1(_00216_),
    .A2(_04843_),
    .B1(_04907_),
    .B2(_00217_),
    .X(_00218_));
 sky130_fd_sc_hd__nand4_1 _07601_ (.A(_00217_),
    .B(_00216_),
    .C(_04843_),
    .D(_04907_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand4_1 _07602_ (.A(_03013_),
    .B(_06613_),
    .C(_00218_),
    .D(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__buf_6 _07603_ (.A(net119),
    .X(_00221_));
 sky130_fd_sc_hd__a22o_1 _07604_ (.A1(_00221_),
    .A2(_06613_),
    .B1(_00218_),
    .B2(_00219_),
    .X(_00222_));
 sky130_fd_sc_hd__nand3_1 _07605_ (.A(_00215_),
    .B(_00220_),
    .C(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__a21o_1 _07606_ (.A1(_00220_),
    .A2(_00222_),
    .B1(_00215_),
    .X(_00224_));
 sky130_fd_sc_hd__nand3_1 _07607_ (.A(_00214_),
    .B(_00223_),
    .C(_00224_),
    .Y(_00225_));
 sky130_fd_sc_hd__a21o_1 _07608_ (.A1(_00223_),
    .A2(_00224_),
    .B1(_00214_),
    .X(_00226_));
 sky130_fd_sc_hd__a21bo_1 _07609_ (.A1(_00116_),
    .A2(_00117_),
    .B1_N(_00115_),
    .X(_00227_));
 sky130_fd_sc_hd__nand3_1 _07610_ (.A(_00225_),
    .B(_00226_),
    .C(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__a21o_1 _07611_ (.A1(_00225_),
    .A2(_00226_),
    .B1(_00227_),
    .X(_00229_));
 sky130_fd_sc_hd__and3_1 _07612_ (.A(net50),
    .B(net51),
    .C(_04509_),
    .X(_00230_));
 sky130_fd_sc_hd__buf_2 _07613_ (.A(net51),
    .X(_00231_));
 sky130_fd_sc_hd__a22o_1 _07614_ (.A1(_00231_),
    .A2(_00083_),
    .B1(_00098_),
    .B2(_03217_),
    .X(_00232_));
 sky130_fd_sc_hd__a21bo_1 _07615_ (.A1(_00093_),
    .A2(_00230_),
    .B1_N(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__nand2_1 _07616_ (.A(_00077_),
    .B(_04369_),
    .Y(_00234_));
 sky130_fd_sc_hd__xor2_2 _07617_ (.A(_00233_),
    .B(_00234_),
    .X(_00235_));
 sky130_fd_sc_hd__and2_1 _07618_ (.A(_03152_),
    .B(_00047_),
    .X(_00236_));
 sky130_fd_sc_hd__clkbuf_4 _07619_ (.A(net118),
    .X(_00237_));
 sky130_fd_sc_hd__a22o_1 _07620_ (.A1(_00081_),
    .A2(_04638_),
    .B1(_04703_),
    .B2(_00237_),
    .X(_00238_));
 sky130_fd_sc_hd__nand4_1 _07621_ (.A(_03056_),
    .B(_03099_),
    .C(_00048_),
    .D(_00033_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand3_1 _07622_ (.A(_00236_),
    .B(_00238_),
    .C(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__a21o_1 _07623_ (.A1(_00238_),
    .A2(_00239_),
    .B1(_00236_),
    .X(_00241_));
 sky130_fd_sc_hd__o21bai_1 _07624_ (.A1(_00131_),
    .A2(_00134_),
    .B1_N(_00130_),
    .Y(_00242_));
 sky130_fd_sc_hd__and3_1 _07625_ (.A(_00240_),
    .B(_00241_),
    .C(_00242_),
    .X(_00243_));
 sky130_fd_sc_hd__a21o_1 _07626_ (.A1(_00240_),
    .A2(_00241_),
    .B1(_00242_),
    .X(_00244_));
 sky130_fd_sc_hd__or2b_1 _07627_ (.A(_00243_),
    .B_N(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__xnor2_2 _07628_ (.A(_00235_),
    .B(_00245_),
    .Y(_00246_));
 sky130_fd_sc_hd__and3_1 _07629_ (.A(_00228_),
    .B(_00229_),
    .C(_00246_),
    .X(_00247_));
 sky130_fd_sc_hd__a21oi_1 _07630_ (.A1(_00228_),
    .A2(_00229_),
    .B1(_00246_),
    .Y(_00248_));
 sky130_fd_sc_hd__a211o_1 _07631_ (.A1(_00020_),
    .A2(_00021_),
    .B1(_00247_),
    .C1(_00248_),
    .X(_00249_));
 sky130_fd_sc_hd__o211ai_1 _07632_ (.A1(_00247_),
    .A2(_00248_),
    .B1(_00020_),
    .C1(_00021_),
    .Y(_00250_));
 sky130_fd_sc_hd__a211o_1 _07633_ (.A1(_00249_),
    .A2(_00250_),
    .B1(_00143_),
    .C1(_00121_),
    .X(_00251_));
 sky130_fd_sc_hd__o211ai_2 _07634_ (.A1(_00121_),
    .A2(_00143_),
    .B1(_00250_),
    .C1(_00249_),
    .Y(_00252_));
 sky130_fd_sc_hd__a22oi_2 _07635_ (.A1(_00212_),
    .A2(_00213_),
    .B1(_00251_),
    .B2(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__and4_1 _07636_ (.A(_00252_),
    .B(_00212_),
    .C(_00213_),
    .D(_00251_),
    .X(_00254_));
 sky130_fd_sc_hd__a211o_2 _07637_ (.A1(_00026_),
    .A2(_00148_),
    .B1(_00253_),
    .C1(_00254_),
    .X(_00255_));
 sky130_fd_sc_hd__o211ai_2 _07638_ (.A1(_00254_),
    .A2(_00253_),
    .B1(_00148_),
    .C1(_00026_),
    .Y(_00256_));
 sky130_fd_sc_hd__and4_1 _07639_ (.A(_00095_),
    .B(_00096_),
    .C(_04358_),
    .D(_04434_),
    .X(_00257_));
 sky130_fd_sc_hd__a22oi_1 _07640_ (.A1(_03099_),
    .A2(_04358_),
    .B1(_04445_),
    .B2(_03056_),
    .Y(_00258_));
 sky130_fd_sc_hd__buf_4 _07641_ (.A(_00074_),
    .X(_00259_));
 sky130_fd_sc_hd__and4bb_1 _07642_ (.A_N(_00257_),
    .B_N(_00258_),
    .C(_03163_),
    .D(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__nor2_1 _07643_ (.A(_00257_),
    .B(_00260_),
    .Y(_00261_));
 sky130_fd_sc_hd__buf_4 _07644_ (.A(_00088_),
    .X(_00262_));
 sky130_fd_sc_hd__o2bb2a_1 _07645_ (.A1_N(_00262_),
    .A2_N(_04369_),
    .B1(_00080_),
    .B2(_00087_),
    .X(_00263_));
 sky130_fd_sc_hd__nor2_1 _07646_ (.A(_00091_),
    .B(_00263_),
    .Y(_00264_));
 sky130_fd_sc_hd__and2b_1 _07647_ (.A_N(_00261_),
    .B(_00264_),
    .X(_00265_));
 sky130_fd_sc_hd__buf_4 _07648_ (.A(net124),
    .X(_00266_));
 sky130_fd_sc_hd__buf_4 _07649_ (.A(_00266_),
    .X(_00267_));
 sky130_fd_sc_hd__and4_1 _07650_ (.A(_03217_),
    .B(_03271_),
    .C(_00267_),
    .D(_04294_),
    .X(_00268_));
 sky130_fd_sc_hd__a22oi_1 _07651_ (.A1(_00125_),
    .A2(_00267_),
    .B1(_04305_),
    .B2(_00124_),
    .Y(_00269_));
 sky130_fd_sc_hd__buf_4 _07652_ (.A(net114),
    .X(_00270_));
 sky130_fd_sc_hd__clkbuf_4 _07653_ (.A(net125),
    .X(_00271_));
 sky130_fd_sc_hd__buf_4 _07654_ (.A(_00271_),
    .X(_00272_));
 sky130_fd_sc_hd__and4bb_1 _07655_ (.A_N(_00268_),
    .B_N(_00269_),
    .C(_00270_),
    .D(_00272_),
    .X(_00273_));
 sky130_fd_sc_hd__o2bb2a_1 _07656_ (.A1_N(_03335_),
    .A2_N(_04186_),
    .B1(_00268_),
    .B2(_00269_),
    .X(_00274_));
 sky130_fd_sc_hd__nor2_1 _07657_ (.A(_00273_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__xnor2_1 _07658_ (.A(_00261_),
    .B(_00264_),
    .Y(_00276_));
 sky130_fd_sc_hd__and2_1 _07659_ (.A(_00275_),
    .B(_00276_),
    .X(_00277_));
 sky130_fd_sc_hd__clkbuf_4 _07660_ (.A(net113),
    .X(_00278_));
 sky130_fd_sc_hd__clkbuf_4 _07661_ (.A(net54),
    .X(_00279_));
 sky130_fd_sc_hd__and4_1 _07662_ (.A(_00278_),
    .B(_00279_),
    .C(_04035_),
    .D(_06433_),
    .X(_00280_));
 sky130_fd_sc_hd__buf_4 _07663_ (.A(net113),
    .X(_00281_));
 sky130_fd_sc_hd__a22oi_1 _07664_ (.A1(_03443_),
    .A2(_06446_),
    .B1(_04111_),
    .B2(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__buf_4 _07665_ (.A(net55),
    .X(_00283_));
 sky130_fd_sc_hd__and4bb_1 _07666_ (.A_N(_00280_),
    .B_N(_00282_),
    .C(_00283_),
    .D(_06437_),
    .X(_00284_));
 sky130_fd_sc_hd__nor2_2 _07667_ (.A(_00280_),
    .B(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__nor2_1 _07668_ (.A(_00268_),
    .B(_00273_),
    .Y(_00286_));
 sky130_fd_sc_hd__clkbuf_4 _07669_ (.A(_04165_),
    .X(_00287_));
 sky130_fd_sc_hd__and4_1 _07670_ (.A(_00278_),
    .B(_03432_),
    .C(_06431_),
    .D(_00287_),
    .X(_00288_));
 sky130_fd_sc_hd__buf_4 _07671_ (.A(_03432_),
    .X(_00289_));
 sky130_fd_sc_hd__buf_4 _07672_ (.A(net113),
    .X(_00290_));
 sky130_fd_sc_hd__a22oi_1 _07673_ (.A1(_00289_),
    .A2(_06433_),
    .B1(_04176_),
    .B2(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__buf_4 _07674_ (.A(net55),
    .X(_00292_));
 sky130_fd_sc_hd__and4bb_1 _07675_ (.A_N(_00288_),
    .B_N(_00291_),
    .C(_00292_),
    .D(_06443_),
    .X(_00293_));
 sky130_fd_sc_hd__o2bb2a_1 _07676_ (.A1_N(_00283_),
    .A2_N(_04046_),
    .B1(_00288_),
    .B2(_00291_),
    .X(_00294_));
 sky130_fd_sc_hd__nor2_1 _07677_ (.A(_00293_),
    .B(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__xnor2_1 _07678_ (.A(_00286_),
    .B(_00295_),
    .Y(_00296_));
 sky130_fd_sc_hd__xnor2_2 _07679_ (.A(_00285_),
    .B(_00296_),
    .Y(_00297_));
 sky130_fd_sc_hd__o21ai_4 _07680_ (.A1(_00265_),
    .A2(_00277_),
    .B1(_00297_),
    .Y(_00298_));
 sky130_fd_sc_hd__buf_2 _07681_ (.A(net50),
    .X(_00299_));
 sky130_fd_sc_hd__and4_1 _07682_ (.A(_00299_),
    .B(_00231_),
    .C(_00287_),
    .D(_00267_),
    .X(_00300_));
 sky130_fd_sc_hd__buf_4 _07683_ (.A(_00267_),
    .X(_00301_));
 sky130_fd_sc_hd__a22oi_1 _07684_ (.A1(_03282_),
    .A2(_04176_),
    .B1(_00301_),
    .B2(_00124_),
    .Y(_00302_));
 sky130_fd_sc_hd__clkbuf_4 _07685_ (.A(_06433_),
    .X(_00303_));
 sky130_fd_sc_hd__and4bb_1 _07686_ (.A_N(_00300_),
    .B_N(_00302_),
    .C(_00270_),
    .D(_00303_),
    .X(_00304_));
 sky130_fd_sc_hd__nor2_1 _07687_ (.A(_00300_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__o2bb2a_1 _07688_ (.A1_N(_00283_),
    .A2_N(_03971_),
    .B1(_00280_),
    .B2(_00282_),
    .X(_00306_));
 sky130_fd_sc_hd__nor2_1 _07689_ (.A(_00284_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__and2b_1 _07690_ (.A_N(_00305_),
    .B(_00307_),
    .X(_00308_));
 sky130_fd_sc_hd__and4_1 _07691_ (.A(_00278_),
    .B(_03432_),
    .C(net132),
    .D(_06430_),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_1 _07692_ (.A(net55),
    .B(net115),
    .Y(_00310_));
 sky130_fd_sc_hd__a22oi_1 _07693_ (.A1(_00279_),
    .A2(_06436_),
    .B1(_04035_),
    .B2(_03378_),
    .Y(_00311_));
 sky130_fd_sc_hd__or3_1 _07694_ (.A(_00309_),
    .B(_00310_),
    .C(_00311_),
    .X(_00312_));
 sky130_fd_sc_hd__and2b_1 _07695_ (.A_N(_00309_),
    .B(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__xnor2_1 _07696_ (.A(_00305_),
    .B(_00307_),
    .Y(_00314_));
 sky130_fd_sc_hd__and2b_1 _07697_ (.A_N(_00313_),
    .B(_00314_),
    .X(_00315_));
 sky130_fd_sc_hd__or3_2 _07698_ (.A(_00265_),
    .B(_00277_),
    .C(_00297_),
    .X(_00316_));
 sky130_fd_sc_hd__o211ai_4 _07699_ (.A1(_00308_),
    .A2(_00315_),
    .B1(_00316_),
    .C1(_00298_),
    .Y(_00317_));
 sky130_fd_sc_hd__and2b_1 _07700_ (.A_N(_00092_),
    .B(_00101_),
    .X(_00318_));
 sky130_fd_sc_hd__or2_1 _07701_ (.A(_00288_),
    .B(_00293_),
    .X(_00319_));
 sky130_fd_sc_hd__nor2_1 _07702_ (.A(_00073_),
    .B(_00076_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(_00292_),
    .B(_04111_),
    .Y(_00321_));
 sky130_fd_sc_hd__and4_1 _07704_ (.A(net113),
    .B(net54),
    .C(_04165_),
    .D(_00266_),
    .X(_00322_));
 sky130_fd_sc_hd__a22o_1 _07705_ (.A1(_03432_),
    .A2(_04165_),
    .B1(_04229_),
    .B2(net113),
    .X(_00323_));
 sky130_fd_sc_hd__and2b_1 _07706_ (.A_N(_00322_),
    .B(_00323_),
    .X(_00324_));
 sky130_fd_sc_hd__xnor2_1 _07707_ (.A(_00321_),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__xnor2_2 _07708_ (.A(_00320_),
    .B(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__xor2_2 _07709_ (.A(_00319_),
    .B(_00326_),
    .X(_00327_));
 sky130_fd_sc_hd__o21ai_2 _07710_ (.A1(_00318_),
    .A2(_00103_),
    .B1(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__or3_1 _07711_ (.A(_00318_),
    .B(_00103_),
    .C(_00327_),
    .X(_00329_));
 sky130_fd_sc_hd__and2b_1 _07712_ (.A_N(_00285_),
    .B(_00296_),
    .X(_00330_));
 sky130_fd_sc_hd__and2b_1 _07713_ (.A_N(_00286_),
    .B(_00295_),
    .X(_00331_));
 sky130_fd_sc_hd__a211oi_2 _07714_ (.A1(_00328_),
    .A2(_00329_),
    .B1(_00330_),
    .C1(_00331_),
    .Y(_00332_));
 sky130_fd_sc_hd__o211a_1 _07715_ (.A1(_00331_),
    .A2(_00330_),
    .B1(_00329_),
    .C1(_00328_),
    .X(_00333_));
 sky130_fd_sc_hd__a211o_1 _07716_ (.A1(_00298_),
    .A2(_00317_),
    .B1(_00332_),
    .C1(_00333_),
    .X(_00334_));
 sky130_fd_sc_hd__a211oi_1 _07717_ (.A1(_00298_),
    .A2(_00317_),
    .B1(_00332_),
    .C1(_00333_),
    .Y(_00335_));
 sky130_fd_sc_hd__o211a_1 _07718_ (.A1(_00333_),
    .A2(_00332_),
    .B1(_00317_),
    .C1(_00298_),
    .X(_00336_));
 sky130_fd_sc_hd__nor2_1 _07719_ (.A(_06455_),
    .B(_06456_),
    .Y(_00337_));
 sky130_fd_sc_hd__or2_1 _07720_ (.A(_06457_),
    .B(_00337_),
    .X(_00338_));
 sky130_fd_sc_hd__or3_2 _07721_ (.A(_00335_),
    .B(_00336_),
    .C(_00338_),
    .X(_00339_));
 sky130_fd_sc_hd__a211oi_1 _07722_ (.A1(_00069_),
    .A2(_00106_),
    .B1(_00144_),
    .C1(_00145_),
    .Y(_00340_));
 sky130_fd_sc_hd__inv_2 _07723_ (.A(_00328_),
    .Y(_00341_));
 sky130_fd_sc_hd__and2b_1 _07724_ (.A_N(_00320_),
    .B(_00325_),
    .X(_00342_));
 sky130_fd_sc_hd__a21oi_2 _07725_ (.A1(_00319_),
    .A2(_00326_),
    .B1(_00342_),
    .Y(_00343_));
 sky130_fd_sc_hd__a32o_1 _07726_ (.A1(_03324_),
    .A2(_04316_),
    .A3(_00127_),
    .B1(_00126_),
    .B2(_04380_),
    .X(_00344_));
 sky130_fd_sc_hd__buf_4 _07727_ (.A(net55),
    .X(_00345_));
 sky130_fd_sc_hd__a22o_1 _07728_ (.A1(_03443_),
    .A2(_04240_),
    .B1(_04305_),
    .B2(_00290_),
    .X(_00346_));
 sky130_fd_sc_hd__nand4_1 _07729_ (.A(_00281_),
    .B(_03443_),
    .C(_04240_),
    .D(_04305_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand4_1 _07730_ (.A(_00345_),
    .B(_04186_),
    .C(_00346_),
    .D(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__a22o_1 _07731_ (.A1(_03486_),
    .A2(_04186_),
    .B1(_00346_),
    .B2(_00347_),
    .X(_00349_));
 sky130_fd_sc_hd__nand3_1 _07732_ (.A(_00344_),
    .B(_00348_),
    .C(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__a31o_1 _07733_ (.A1(_03497_),
    .A2(_04122_),
    .A3(_00323_),
    .B1(_00322_),
    .X(_00351_));
 sky130_fd_sc_hd__a21o_1 _07734_ (.A1(_00348_),
    .A2(_00349_),
    .B1(_00344_),
    .X(_00352_));
 sky130_fd_sc_hd__nand3_1 _07735_ (.A(_00350_),
    .B(_00351_),
    .C(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__a21o_1 _07736_ (.A1(_00129_),
    .A2(_00139_),
    .B1(_00138_),
    .X(_00354_));
 sky130_fd_sc_hd__a21o_1 _07737_ (.A1(_00350_),
    .A2(_00352_),
    .B1(_00351_),
    .X(_00355_));
 sky130_fd_sc_hd__and3_1 _07738_ (.A(_00353_),
    .B(_00354_),
    .C(_00355_),
    .X(_00356_));
 sky130_fd_sc_hd__a21oi_1 _07739_ (.A1(_00353_),
    .A2(_00355_),
    .B1(_00354_),
    .Y(_00357_));
 sky130_fd_sc_hd__nor2_1 _07740_ (.A(_00356_),
    .B(_00357_),
    .Y(_00358_));
 sky130_fd_sc_hd__xnor2_2 _07741_ (.A(_00343_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__o21a_1 _07742_ (.A1(_00341_),
    .A2(_00333_),
    .B1(_00359_),
    .X(_00360_));
 sky130_fd_sc_hd__nor3_1 _07743_ (.A(_00341_),
    .B(_00333_),
    .C(_00359_),
    .Y(_00361_));
 sky130_fd_sc_hd__nor2_1 _07744_ (.A(_06452_),
    .B(_06457_),
    .Y(_00362_));
 sky130_fd_sc_hd__or2_1 _07745_ (.A(_06458_),
    .B(_00362_),
    .X(_00363_));
 sky130_fd_sc_hd__o21ai_1 _07746_ (.A1(_00360_),
    .A2(_00361_),
    .B1(_00363_),
    .Y(_00364_));
 sky130_fd_sc_hd__or3_1 _07747_ (.A(_00360_),
    .B(_00361_),
    .C(_00363_),
    .X(_00365_));
 sky130_fd_sc_hd__o211a_1 _07748_ (.A1(_00144_),
    .A2(_00340_),
    .B1(_00364_),
    .C1(_00365_),
    .X(_00366_));
 sky130_fd_sc_hd__a211oi_1 _07749_ (.A1(_00365_),
    .A2(_00364_),
    .B1(_00340_),
    .C1(_00144_),
    .Y(_00367_));
 sky130_fd_sc_hd__a211o_1 _07750_ (.A1(_00334_),
    .A2(_00339_),
    .B1(_00366_),
    .C1(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__o211ai_2 _07751_ (.A1(_00366_),
    .A2(_00367_),
    .B1(_00334_),
    .C1(_00339_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand4_2 _07752_ (.A(_00255_),
    .B(_00256_),
    .C(_00368_),
    .D(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand4_1 _07753_ (.A(_00252_),
    .B(_00212_),
    .C(_00213_),
    .D(_00251_),
    .Y(_00371_));
 sky130_fd_sc_hd__nor3_1 _07754_ (.A(_00186_),
    .B(_00187_),
    .C(_00209_),
    .Y(_00372_));
 sky130_fd_sc_hd__and3_1 _07755_ (.A(_00168_),
    .B(_00169_),
    .C(_00170_),
    .X(_00373_));
 sky130_fd_sc_hd__nand4_1 _07756_ (.A(_06534_),
    .B(_02205_),
    .C(_00153_),
    .D(net29),
    .Y(_00374_));
 sky130_fd_sc_hd__and2_1 _07757_ (.A(_06460_),
    .B(net128),
    .X(_00375_));
 sky130_fd_sc_hd__a22o_1 _07758_ (.A1(_02205_),
    .A2(_00153_),
    .B1(net29),
    .B2(_06534_),
    .X(_00376_));
 sky130_fd_sc_hd__nand3_1 _07759_ (.A(_00374_),
    .B(_00375_),
    .C(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__o21bai_1 _07760_ (.A1(_00152_),
    .A2(_00154_),
    .B1_N(_00151_),
    .Y(_00378_));
 sky130_fd_sc_hd__a21o_1 _07761_ (.A1(_00374_),
    .A2(_00376_),
    .B1(_00375_),
    .X(_00379_));
 sky130_fd_sc_hd__nand3_1 _07762_ (.A(_00377_),
    .B(_00378_),
    .C(_00379_),
    .Y(_00380_));
 sky130_fd_sc_hd__a21o_1 _07763_ (.A1(_00377_),
    .A2(_00379_),
    .B1(_00378_),
    .X(_00381_));
 sky130_fd_sc_hd__clkbuf_4 _07764_ (.A(_05627_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(_06544_),
    .B(_00382_),
    .Y(_00383_));
 sky130_fd_sc_hd__and4_1 _07766_ (.A(_06503_),
    .B(_06504_),
    .C(net130),
    .D(net129),
    .X(_00384_));
 sky130_fd_sc_hd__clkbuf_4 _07767_ (.A(net129),
    .X(_00385_));
 sky130_fd_sc_hd__a22oi_1 _07768_ (.A1(_00162_),
    .A2(_00163_),
    .B1(_00385_),
    .B2(_00164_),
    .Y(_00386_));
 sky130_fd_sc_hd__nor2_1 _07769_ (.A(_00384_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_00383_),
    .B(_00387_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand3_1 _07771_ (.A(_00380_),
    .B(_00381_),
    .C(_00388_),
    .Y(_00389_));
 sky130_fd_sc_hd__a21bo_1 _07772_ (.A1(_00159_),
    .A2(_00167_),
    .B1_N(_00158_),
    .X(_00390_));
 sky130_fd_sc_hd__a21o_1 _07773_ (.A1(_00380_),
    .A2(_00381_),
    .B1(_00388_),
    .X(_00391_));
 sky130_fd_sc_hd__nand3_1 _07774_ (.A(_00389_),
    .B(_00390_),
    .C(_00391_),
    .Y(_00392_));
 sky130_fd_sc_hd__a21o_1 _07775_ (.A1(_00389_),
    .A2(_00391_),
    .B1(_00390_),
    .X(_00393_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(_00177_),
    .B(_00178_),
    .Y(_00394_));
 sky130_fd_sc_hd__o21bai_1 _07777_ (.A1(_00160_),
    .A2(_00165_),
    .B1_N(_00161_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _07778_ (.A(_06663_),
    .B(_06666_),
    .Y(_00396_));
 sky130_fd_sc_hd__a22o_1 _07779_ (.A1(_06516_),
    .A2(_05498_),
    .B1(_05563_),
    .B2(_06520_),
    .X(_00397_));
 sky130_fd_sc_hd__buf_4 _07780_ (.A(_06466_),
    .X(_00398_));
 sky130_fd_sc_hd__nand4_1 _07781_ (.A(_06565_),
    .B(_02485_),
    .C(_00398_),
    .D(_05563_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand3b_1 _07782_ (.A_N(_00396_),
    .B(_00397_),
    .C(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__a21bo_1 _07783_ (.A1(_00397_),
    .A2(_00399_),
    .B1_N(_00396_),
    .X(_00401_));
 sky130_fd_sc_hd__and3_1 _07784_ (.A(_00395_),
    .B(_00400_),
    .C(_00401_),
    .X(_00402_));
 sky130_fd_sc_hd__a21o_1 _07785_ (.A1(_00400_),
    .A2(_00401_),
    .B1(_00395_),
    .X(_00403_));
 sky130_fd_sc_hd__and2b_1 _07786_ (.A_N(_00402_),
    .B(_00403_),
    .X(_00404_));
 sky130_fd_sc_hd__xor2_1 _07787_ (.A(_00394_),
    .B(_00404_),
    .X(_00405_));
 sky130_fd_sc_hd__a21o_1 _07788_ (.A1(_00392_),
    .A2(_00393_),
    .B1(_00405_),
    .X(_00406_));
 sky130_fd_sc_hd__nand3_1 _07789_ (.A(_00392_),
    .B(_00393_),
    .C(_00405_),
    .Y(_00407_));
 sky130_fd_sc_hd__o211ai_2 _07790_ (.A1(_00373_),
    .A2(_00185_),
    .B1(_00406_),
    .C1(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__a211o_1 _07791_ (.A1(_00407_),
    .A2(_00406_),
    .B1(_00185_),
    .C1(_00373_),
    .X(_00409_));
 sky130_fd_sc_hd__a21o_1 _07792_ (.A1(_00173_),
    .A2(_00181_),
    .B1(_00180_),
    .X(_00410_));
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(_02712_),
    .B(_06568_),
    .Y(_00411_));
 sky130_fd_sc_hd__buf_4 _07794_ (.A(_05305_),
    .X(_00412_));
 sky130_fd_sc_hd__a22oi_2 _07795_ (.A1(_06682_),
    .A2(_00412_),
    .B1(_05380_),
    .B2(_00000_),
    .Y(_00413_));
 sky130_fd_sc_hd__buf_6 _07796_ (.A(net68),
    .X(_00414_));
 sky130_fd_sc_hd__and4_1 _07797_ (.A(_00414_),
    .B(_06622_),
    .C(_05305_),
    .D(_05370_),
    .X(_00415_));
 sky130_fd_sc_hd__or3_1 _07798_ (.A(_00411_),
    .B(_00413_),
    .C(_00415_),
    .X(_00416_));
 sky130_fd_sc_hd__o21ai_1 _07799_ (.A1(_00413_),
    .A2(_00415_),
    .B1(_00411_),
    .Y(_00417_));
 sky130_fd_sc_hd__o21bai_1 _07800_ (.A1(_00189_),
    .A2(_00190_),
    .B1_N(_00191_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand3_1 _07801_ (.A(_00416_),
    .B(_00417_),
    .C(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(_00416_),
    .A2(_00417_),
    .B1(_00418_),
    .X(_00420_));
 sky130_fd_sc_hd__buf_4 _07803_ (.A(_06584_),
    .X(_00421_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(_02840_),
    .B(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__buf_4 _07805_ (.A(_05112_),
    .X(_00423_));
 sky130_fd_sc_hd__a22oi_2 _07806_ (.A1(_02808_),
    .A2(_00423_),
    .B1(_00002_),
    .B2(_02765_),
    .Y(_00424_));
 sky130_fd_sc_hd__and4_1 _07807_ (.A(_06606_),
    .B(_06601_),
    .C(_05112_),
    .D(_05187_),
    .X(_00425_));
 sky130_fd_sc_hd__nor2_1 _07808_ (.A(_00424_),
    .B(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__xnor2_1 _07809_ (.A(_00422_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand3_1 _07810_ (.A(_00419_),
    .B(_00420_),
    .C(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__a21o_1 _07811_ (.A1(_00419_),
    .A2(_00420_),
    .B1(_00427_),
    .X(_00429_));
 sky130_fd_sc_hd__nand3_1 _07812_ (.A(_00410_),
    .B(_00428_),
    .C(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(_00195_),
    .B(_00202_),
    .Y(_00431_));
 sky130_fd_sc_hd__a21o_1 _07814_ (.A1(_00428_),
    .A2(_00429_),
    .B1(_00410_),
    .X(_00432_));
 sky130_fd_sc_hd__nand3_1 _07815_ (.A(_00430_),
    .B(_00431_),
    .C(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__a21o_1 _07816_ (.A1(_00430_),
    .A2(_00432_),
    .B1(_00431_),
    .X(_00434_));
 sky130_fd_sc_hd__and2_1 _07817_ (.A(_00433_),
    .B(_00434_),
    .X(_00435_));
 sky130_fd_sc_hd__a21o_1 _07818_ (.A1(_00408_),
    .A2(_00409_),
    .B1(_00435_),
    .X(_00436_));
 sky130_fd_sc_hd__nand3_1 _07819_ (.A(_00408_),
    .B(_00409_),
    .C(_00435_),
    .Y(_00437_));
 sky130_fd_sc_hd__o211ai_1 _07820_ (.A1(_00186_),
    .A2(_00372_),
    .B1(_00436_),
    .C1(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__a211o_1 _07821_ (.A1(_00437_),
    .A2(_00436_),
    .B1(_00372_),
    .C1(_00186_),
    .X(_00439_));
 sky130_fd_sc_hd__inv_2 _07822_ (.A(_00228_),
    .Y(_00440_));
 sky130_fd_sc_hd__nor2_1 _07823_ (.A(_00440_),
    .B(_00247_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _07824_ (.A(_00219_),
    .B(_00220_),
    .Y(_00442_));
 sky130_fd_sc_hd__a32o_1 _07825_ (.A1(_02840_),
    .A2(_00197_),
    .A3(_00199_),
    .B1(_00010_),
    .B2(_05123_),
    .X(_00443_));
 sky130_fd_sc_hd__buf_6 _07826_ (.A(net45),
    .X(_00444_));
 sky130_fd_sc_hd__buf_6 _07827_ (.A(_06603_),
    .X(_00445_));
 sky130_fd_sc_hd__a22o_1 _07828_ (.A1(_00046_),
    .A2(_06605_),
    .B1(_06591_),
    .B2(_00049_),
    .X(_00446_));
 sky130_fd_sc_hd__nand4_1 _07829_ (.A(_00063_),
    .B(_00216_),
    .C(_06605_),
    .D(_06591_),
    .Y(_00447_));
 sky130_fd_sc_hd__a22o_1 _07830_ (.A1(_00444_),
    .A2(_00445_),
    .B1(_00446_),
    .B2(_00447_),
    .X(_00448_));
 sky130_fd_sc_hd__nand4_1 _07831_ (.A(_00221_),
    .B(_04854_),
    .C(_00446_),
    .D(_00447_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand3_1 _07832_ (.A(_00443_),
    .B(_00448_),
    .C(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__a21o_1 _07833_ (.A1(_00448_),
    .A2(_00449_),
    .B1(_00443_),
    .X(_00451_));
 sky130_fd_sc_hd__nand3_1 _07834_ (.A(_00442_),
    .B(_00450_),
    .C(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__a21o_1 _07835_ (.A1(_00450_),
    .A2(_00451_),
    .B1(_00442_),
    .X(_00453_));
 sky130_fd_sc_hd__a21bo_1 _07836_ (.A1(_00214_),
    .A2(_00224_),
    .B1_N(_00223_),
    .X(_00454_));
 sky130_fd_sc_hd__and3_1 _07837_ (.A(_00452_),
    .B(_00453_),
    .C(_00454_),
    .X(_00455_));
 sky130_fd_sc_hd__a21oi_1 _07838_ (.A1(_00452_),
    .A2(_00453_),
    .B1(_00454_),
    .Y(_00456_));
 sky130_fd_sc_hd__a22o_1 _07839_ (.A1(_03271_),
    .A2(_04509_),
    .B1(_00035_),
    .B2(_03217_),
    .X(_00457_));
 sky130_fd_sc_hd__a21bo_1 _07840_ (.A1(_00036_),
    .A2(_00230_),
    .B1_N(_00457_),
    .X(_00458_));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(_03324_),
    .B(_04456_),
    .Y(_00459_));
 sky130_fd_sc_hd__xor2_2 _07842_ (.A(_00458_),
    .B(_00459_),
    .X(_00460_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_03152_),
    .B(_04638_),
    .Y(_00461_));
 sky130_fd_sc_hd__buf_4 _07844_ (.A(net117),
    .X(_00462_));
 sky130_fd_sc_hd__a22oi_2 _07845_ (.A1(_00462_),
    .A2(_04703_),
    .B1(_04778_),
    .B2(_00237_),
    .Y(_00463_));
 sky130_fd_sc_hd__and4_1 _07846_ (.A(_00095_),
    .B(_00096_),
    .C(_04703_),
    .D(_06611_),
    .X(_00464_));
 sky130_fd_sc_hd__or3_1 _07847_ (.A(_00461_),
    .B(_00463_),
    .C(_00464_),
    .X(_00465_));
 sky130_fd_sc_hd__o21ai_1 _07848_ (.A1(_00463_),
    .A2(_00464_),
    .B1(_00461_),
    .Y(_00466_));
 sky130_fd_sc_hd__a21bo_1 _07849_ (.A1(_00236_),
    .A2(_00238_),
    .B1_N(_00239_),
    .X(_00467_));
 sky130_fd_sc_hd__and3_1 _07850_ (.A(_00465_),
    .B(_00466_),
    .C(_00467_),
    .X(_00468_));
 sky130_fd_sc_hd__a21o_1 _07851_ (.A1(_00465_),
    .A2(_00466_),
    .B1(_00467_),
    .X(_00469_));
 sky130_fd_sc_hd__and2b_1 _07852_ (.A_N(_00468_),
    .B(_00469_),
    .X(_00470_));
 sky130_fd_sc_hd__xnor2_2 _07853_ (.A(_00460_),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__nor3_1 _07854_ (.A(_00455_),
    .B(_00456_),
    .C(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__o21a_1 _07855_ (.A1(_00455_),
    .A2(_00456_),
    .B1(_00471_),
    .X(_00473_));
 sky130_fd_sc_hd__a211oi_1 _07856_ (.A1(_00204_),
    .A2(_00207_),
    .B1(_00472_),
    .C1(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__o211a_1 _07857_ (.A1(_00472_),
    .A2(_00473_),
    .B1(_00204_),
    .C1(_00207_),
    .X(_00475_));
 sky130_fd_sc_hd__nor2_1 _07858_ (.A(_00474_),
    .B(_00475_),
    .Y(_00476_));
 sky130_fd_sc_hd__xnor2_1 _07859_ (.A(_00441_),
    .B(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__a21oi_1 _07860_ (.A1(_00438_),
    .A2(_00439_),
    .B1(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__and3_1 _07861_ (.A(_00438_),
    .B(_00439_),
    .C(_00477_),
    .X(_00479_));
 sky130_fd_sc_hd__a211o_1 _07862_ (.A1(_00212_),
    .A2(_00371_),
    .B1(_00478_),
    .C1(_00479_),
    .X(_00480_));
 sky130_fd_sc_hd__o211ai_2 _07863_ (.A1(_00479_),
    .A2(_00478_),
    .B1(_00371_),
    .C1(_00212_),
    .Y(_00481_));
 sky130_fd_sc_hd__or2b_1 _07864_ (.A(_00360_),
    .B_N(_00365_),
    .X(_00482_));
 sky130_fd_sc_hd__nand2_1 _07865_ (.A(_00249_),
    .B(_00252_),
    .Y(_00483_));
 sky130_fd_sc_hd__a21o_1 _07866_ (.A1(_00235_),
    .A2(_00244_),
    .B1(_00243_),
    .X(_00484_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(_00347_),
    .B(_00348_),
    .Y(_00485_));
 sky130_fd_sc_hd__a32o_1 _07868_ (.A1(_00270_),
    .A2(_04369_),
    .A3(_00232_),
    .B1(_00230_),
    .B2(_04456_),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _07869_ (.A1(_00279_),
    .A2(_00074_),
    .B1(_00090_),
    .B2(_00278_),
    .X(_00487_));
 sky130_fd_sc_hd__nand4_2 _07870_ (.A(_03378_),
    .B(_00289_),
    .C(_00074_),
    .D(_00090_),
    .Y(_00488_));
 sky130_fd_sc_hd__a22o_1 _07871_ (.A1(_00292_),
    .A2(_00301_),
    .B1(_00487_),
    .B2(_00488_),
    .X(_00489_));
 sky130_fd_sc_hd__nand4_2 _07872_ (.A(_00283_),
    .B(_04251_),
    .C(_00487_),
    .D(_00488_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand3_2 _07873_ (.A(_00486_),
    .B(_00489_),
    .C(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__a21o_1 _07874_ (.A1(_00489_),
    .A2(_00490_),
    .B1(_00486_),
    .X(_00492_));
 sky130_fd_sc_hd__nand3_1 _07875_ (.A(_00485_),
    .B(_00491_),
    .C(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__a21o_1 _07876_ (.A1(_00491_),
    .A2(_00492_),
    .B1(_00485_),
    .X(_00494_));
 sky130_fd_sc_hd__and3_1 _07877_ (.A(_00484_),
    .B(_00493_),
    .C(_00494_),
    .X(_00495_));
 sky130_fd_sc_hd__a21oi_1 _07878_ (.A1(_00493_),
    .A2(_00494_),
    .B1(_00484_),
    .Y(_00496_));
 sky130_fd_sc_hd__a211oi_1 _07879_ (.A1(_00350_),
    .A2(_00353_),
    .B1(_00495_),
    .C1(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__o211a_1 _07880_ (.A1(_00495_),
    .A2(_00496_),
    .B1(_00350_),
    .C1(_00353_),
    .X(_00498_));
 sky130_fd_sc_hd__or2_1 _07881_ (.A(_00497_),
    .B(_00498_),
    .X(_00499_));
 sky130_fd_sc_hd__o21ba_1 _07882_ (.A1(_00343_),
    .A2(_00357_),
    .B1_N(_00356_),
    .X(_00500_));
 sky130_fd_sc_hd__xnor2_2 _07883_ (.A(_00499_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__clkbuf_4 _07884_ (.A(net61),
    .X(_00502_));
 sky130_fd_sc_hd__nand2_2 _07885_ (.A(_00502_),
    .B(_03917_),
    .Y(_00503_));
 sky130_fd_sc_hd__and2_1 _07886_ (.A(_06441_),
    .B(_06448_),
    .X(_00504_));
 sky130_fd_sc_hd__nand2_1 _07887_ (.A(_03722_),
    .B(_03993_),
    .Y(_00505_));
 sky130_fd_sc_hd__buf_2 _07888_ (.A(net112),
    .X(_00506_));
 sky130_fd_sc_hd__a22oi_1 _07889_ (.A1(_03604_),
    .A2(_06433_),
    .B1(_00272_),
    .B2(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__and4_1 _07890_ (.A(net112),
    .B(_03593_),
    .C(_06431_),
    .D(_00287_),
    .X(_00508_));
 sky130_fd_sc_hd__and4bb_1 _07891_ (.A_N(_00507_),
    .B_N(_00508_),
    .C(_06439_),
    .D(_06443_),
    .X(_00509_));
 sky130_fd_sc_hd__o2bb2a_1 _07892_ (.A1_N(_06439_),
    .A2_N(_04046_),
    .B1(_00507_),
    .B2(_00508_),
    .X(_00510_));
 sky130_fd_sc_hd__nor2_1 _07893_ (.A(_00509_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__nor2_1 _07894_ (.A(_06432_),
    .B(_06438_),
    .Y(_00512_));
 sky130_fd_sc_hd__xnor2_1 _07895_ (.A(_00511_),
    .B(_00512_),
    .Y(_00513_));
 sky130_fd_sc_hd__xnor2_1 _07896_ (.A(_00505_),
    .B(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__o21a_1 _07897_ (.A1(_00504_),
    .A2(_06450_),
    .B1(_00514_),
    .X(_00515_));
 sky130_fd_sc_hd__or3_1 _07898_ (.A(_00514_),
    .B(_00504_),
    .C(_06450_),
    .X(_00516_));
 sky130_fd_sc_hd__and2b_1 _07899_ (.A_N(_00515_),
    .B(_00516_),
    .X(_00517_));
 sky130_fd_sc_hd__xnor2_4 _07900_ (.A(_00503_),
    .B(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__xnor2_4 _07901_ (.A(_00501_),
    .B(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__xnor2_1 _07902_ (.A(_00483_),
    .B(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__xnor2_2 _07903_ (.A(_00482_),
    .B(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__a21oi_2 _07904_ (.A1(_00480_),
    .A2(_00481_),
    .B1(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__and3_1 _07905_ (.A(_00480_),
    .B(_00481_),
    .C(_00521_),
    .X(_00523_));
 sky130_fd_sc_hd__a211o_1 _07906_ (.A1(_00255_),
    .A2(_00370_),
    .B1(_00522_),
    .C1(_00523_),
    .X(_00524_));
 sky130_fd_sc_hd__or2b_1 _07907_ (.A(_00366_),
    .B_N(_00368_),
    .X(_00525_));
 sky130_fd_sc_hd__o211ai_4 _07908_ (.A1(_00523_),
    .A2(_00522_),
    .B1(_00370_),
    .C1(_00255_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand3_1 _07909_ (.A(_00524_),
    .B(_00525_),
    .C(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__a21o_1 _07910_ (.A1(_00524_),
    .A2(_00526_),
    .B1(_00525_),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _07911_ (.A(_02377_),
    .B(_06561_),
    .Y(_00529_));
 sky130_fd_sc_hd__buf_4 _07912_ (.A(_05370_),
    .X(_00530_));
 sky130_fd_sc_hd__a22oi_2 _07913_ (.A1(_00162_),
    .A2(_00412_),
    .B1(_00530_),
    .B2(_00164_),
    .Y(_00531_));
 sky130_fd_sc_hd__and4_1 _07914_ (.A(_06501_),
    .B(_06500_),
    .C(_06562_),
    .D(_05370_),
    .X(_00532_));
 sky130_fd_sc_hd__o21ba_1 _07915_ (.A1(_00529_),
    .A2(_00531_),
    .B1_N(_00532_),
    .X(_00533_));
 sky130_fd_sc_hd__clkbuf_8 _07916_ (.A(_06623_),
    .X(_00534_));
 sky130_fd_sc_hd__o2bb2a_1 _07917_ (.A1_N(_02528_),
    .A2_N(_00534_),
    .B1(_06514_),
    .B2(_06521_),
    .X(_00535_));
 sky130_fd_sc_hd__or3_1 _07918_ (.A(_06522_),
    .B(_00533_),
    .C(_00535_),
    .X(_00536_));
 sky130_fd_sc_hd__and4_1 _07919_ (.A(_06564_),
    .B(_02474_),
    .C(_05101_),
    .D(_05176_),
    .X(_00537_));
 sky130_fd_sc_hd__a22oi_1 _07920_ (.A1(_06516_),
    .A2(_05101_),
    .B1(_06517_),
    .B2(_06520_),
    .Y(_00538_));
 sky130_fd_sc_hd__and4bb_1 _07921_ (.A_N(_00537_),
    .B_N(_00538_),
    .C(_06663_),
    .D(_06584_),
    .X(_00539_));
 sky130_fd_sc_hd__nor2_1 _07922_ (.A(_00537_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__nor2_1 _07923_ (.A(_06522_),
    .B(_00535_),
    .Y(_00541_));
 sky130_fd_sc_hd__xnor2_1 _07924_ (.A(_00533_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__or2b_1 _07925_ (.A(_00540_),
    .B_N(_00542_),
    .X(_00543_));
 sky130_fd_sc_hd__xnor2_1 _07926_ (.A(_06597_),
    .B(_06615_),
    .Y(_00544_));
 sky130_fd_sc_hd__a21o_2 _07927_ (.A1(_00536_),
    .A2(_00543_),
    .B1(_00544_),
    .X(_00545_));
 sky130_fd_sc_hd__and4_1 _07928_ (.A(_00414_),
    .B(_06579_),
    .C(_04896_),
    .D(_06580_),
    .X(_00546_));
 sky130_fd_sc_hd__a22oi_1 _07929_ (.A1(_02658_),
    .A2(_04896_),
    .B1(_04961_),
    .B2(_02593_),
    .Y(_00547_));
 sky130_fd_sc_hd__and4bb_1 _07930_ (.A_N(_00546_),
    .B_N(_00547_),
    .C(_06593_),
    .D(_04843_),
    .X(_00548_));
 sky130_fd_sc_hd__nor2_1 _07931_ (.A(_00546_),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__buf_4 _07932_ (.A(_04896_),
    .X(_00550_));
 sky130_fd_sc_hd__o2bb2a_1 _07933_ (.A1_N(_06620_),
    .A2_N(_00550_),
    .B1(_06582_),
    .B2(_06586_),
    .X(_00551_));
 sky130_fd_sc_hd__nor2_1 _07934_ (.A(_06587_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__and2b_1 _07935_ (.A_N(_00549_),
    .B(_00552_),
    .X(_00553_));
 sky130_fd_sc_hd__xnor2_1 _07936_ (.A(_00549_),
    .B(_00552_),
    .Y(_00554_));
 sky130_fd_sc_hd__and2_4 _07937_ (.A(_00011_),
    .B(_06612_),
    .X(_00555_));
 sky130_fd_sc_hd__a21oi_1 _07938_ (.A1(_02765_),
    .A2(_04854_),
    .B1(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__o2bb2a_1 _07939_ (.A1_N(_06610_),
    .A2_N(_04725_),
    .B1(_00038_),
    .B2(_00556_),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(_00041_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__and2_1 _07941_ (.A(_00554_),
    .B(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__nand3_1 _07942_ (.A(_00536_),
    .B(_00543_),
    .C(_00544_),
    .Y(_00560_));
 sky130_fd_sc_hd__o211ai_4 _07943_ (.A1(_00553_),
    .A2(_00559_),
    .B1(_00545_),
    .C1(_00560_),
    .Y(_00561_));
 sky130_fd_sc_hd__o21a_1 _07944_ (.A1(_00070_),
    .A2(_00071_),
    .B1(_00105_),
    .X(_00562_));
 sky130_fd_sc_hd__nor3_2 _07945_ (.A(_00070_),
    .B(_00071_),
    .C(_00105_),
    .Y(_00563_));
 sky130_fd_sc_hd__a211oi_4 _07946_ (.A1(_00545_),
    .A2(_00561_),
    .B1(_00562_),
    .C1(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hd__a22o_1 _07947_ (.A1(_00011_),
    .A2(_00040_),
    .B1(_04789_),
    .B2(_00012_),
    .X(_00565_));
 sky130_fd_sc_hd__and2_4 _07948_ (.A(_00012_),
    .B(_00040_),
    .X(_00566_));
 sky130_fd_sc_hd__a32o_2 _07949_ (.A1(_02840_),
    .A2(_00059_),
    .A3(_00565_),
    .B1(_00566_),
    .B2(_00555_),
    .X(_00567_));
 sky130_fd_sc_hd__o2bb2a_1 _07950_ (.A1_N(_03002_),
    .A2_N(_04520_),
    .B1(_00045_),
    .B2(_00050_),
    .X(_00568_));
 sky130_fd_sc_hd__nor2_1 _07951_ (.A(_00051_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_00567_),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__and4_1 _07953_ (.A(_02894_),
    .B(_02948_),
    .C(_00098_),
    .D(_00047_),
    .X(_00571_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_03002_),
    .B(_00093_),
    .Y(_00572_));
 sky130_fd_sc_hd__a22oi_2 _07955_ (.A1(_00062_),
    .A2(_00085_),
    .B1(_04585_),
    .B2(_00063_),
    .Y(_00573_));
 sky130_fd_sc_hd__or3_1 _07956_ (.A(_00571_),
    .B(_00572_),
    .C(_00573_),
    .X(_00574_));
 sky130_fd_sc_hd__or2b_1 _07957_ (.A(_00571_),
    .B_N(_00574_),
    .X(_00575_));
 sky130_fd_sc_hd__xor2_1 _07958_ (.A(_00567_),
    .B(_00569_),
    .X(_00576_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(_00575_),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__xnor2_1 _07960_ (.A(_00052_),
    .B(_00054_),
    .Y(_00578_));
 sky130_fd_sc_hd__a21o_1 _07961_ (.A1(_00570_),
    .A2(_00577_),
    .B1(_00578_),
    .X(_00579_));
 sky130_fd_sc_hd__a21oi_1 _07962_ (.A1(_00570_),
    .A2(_00577_),
    .B1(_00578_),
    .Y(_00580_));
 sky130_fd_sc_hd__and3_1 _07963_ (.A(_00570_),
    .B(_00577_),
    .C(_00578_),
    .X(_00581_));
 sky130_fd_sc_hd__nor2_1 _07964_ (.A(_00275_),
    .B(_00276_),
    .Y(_00582_));
 sky130_fd_sc_hd__or2_1 _07965_ (.A(_00277_),
    .B(_00582_),
    .X(_00583_));
 sky130_fd_sc_hd__or3_1 _07966_ (.A(_00580_),
    .B(_00581_),
    .C(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__o211a_1 _07967_ (.A1(_00563_),
    .A2(_00562_),
    .B1(_00561_),
    .C1(_00545_),
    .X(_00585_));
 sky130_fd_sc_hd__a211oi_1 _07968_ (.A1(_00579_),
    .A2(_00584_),
    .B1(_00564_),
    .C1(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__o21ai_1 _07969_ (.A1(_00335_),
    .A2(_00336_),
    .B1(_00338_),
    .Y(_00587_));
 sky130_fd_sc_hd__o211a_1 _07970_ (.A1(_00564_),
    .A2(_00586_),
    .B1(_00587_),
    .C1(_00339_),
    .X(_00588_));
 sky130_fd_sc_hd__o2bb2a_1 _07971_ (.A1_N(_03335_),
    .A2_N(_04122_),
    .B1(_00300_),
    .B2(_00302_),
    .X(_00589_));
 sky130_fd_sc_hd__nor2_1 _07972_ (.A(_00304_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__o2bb2a_1 _07973_ (.A1_N(_00262_),
    .A2_N(_04316_),
    .B1(_00257_),
    .B2(_00258_),
    .X(_00591_));
 sky130_fd_sc_hd__buf_4 _07974_ (.A(net123),
    .X(_00592_));
 sky130_fd_sc_hd__and4_1 _07975_ (.A(net118),
    .B(net117),
    .C(_00592_),
    .D(_00089_),
    .X(_00593_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_03152_),
    .B(_00267_),
    .Y(_00594_));
 sky130_fd_sc_hd__a22oi_2 _07977_ (.A1(_00096_),
    .A2(_04294_),
    .B1(_04358_),
    .B2(_00095_),
    .Y(_00595_));
 sky130_fd_sc_hd__or3_2 _07978_ (.A(_00593_),
    .B(_00594_),
    .C(_00595_),
    .X(_00596_));
 sky130_fd_sc_hd__and2b_1 _07979_ (.A_N(_00593_),
    .B(_00596_),
    .X(_00597_));
 sky130_fd_sc_hd__o21ai_1 _07980_ (.A1(_00260_),
    .A2(_00591_),
    .B1(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__or3_1 _07981_ (.A(_00260_),
    .B(_00597_),
    .C(_00591_),
    .X(_00599_));
 sky130_fd_sc_hd__a21boi_2 _07982_ (.A1(_00590_),
    .A2(_00598_),
    .B1_N(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__xnor2_1 _07983_ (.A(_00313_),
    .B(_00314_),
    .Y(_00601_));
 sky130_fd_sc_hd__and2b_1 _07984_ (.A_N(_00600_),
    .B(_00601_),
    .X(_00602_));
 sky130_fd_sc_hd__o21ai_1 _07985_ (.A1(_00309_),
    .A2(_00311_),
    .B1(_00310_),
    .Y(_00603_));
 sky130_fd_sc_hd__a22o_1 _07986_ (.A1(_00125_),
    .A2(_06433_),
    .B1(_04176_),
    .B2(_00299_),
    .X(_00604_));
 sky130_fd_sc_hd__and4_1 _07987_ (.A(_00299_),
    .B(_00231_),
    .C(_06433_),
    .D(_00287_),
    .X(_00605_));
 sky130_fd_sc_hd__a31o_1 _07988_ (.A1(_03324_),
    .A2(_04046_),
    .A3(_00604_),
    .B1(_00605_),
    .X(_00606_));
 sky130_fd_sc_hd__a21o_1 _07989_ (.A1(_00312_),
    .A2(_00603_),
    .B1(_00606_),
    .X(_00607_));
 sky130_fd_sc_hd__and4_1 _07990_ (.A(_03389_),
    .B(_03454_),
    .C(_03873_),
    .D(_03971_),
    .X(_00608_));
 sky130_fd_sc_hd__and3_1 _07991_ (.A(_00312_),
    .B(_00606_),
    .C(_00603_),
    .X(_00609_));
 sky130_fd_sc_hd__a21o_1 _07992_ (.A1(_00607_),
    .A2(_00608_),
    .B1(_00609_),
    .X(_00610_));
 sky130_fd_sc_hd__xnor2_1 _07993_ (.A(_00600_),
    .B(_00601_),
    .Y(_00611_));
 sky130_fd_sc_hd__and2_1 _07994_ (.A(_00610_),
    .B(_00611_),
    .X(_00612_));
 sky130_fd_sc_hd__a211o_1 _07995_ (.A1(_00298_),
    .A2(_00316_),
    .B1(_00315_),
    .C1(_00308_),
    .X(_00613_));
 sky130_fd_sc_hd__o211ai_4 _07996_ (.A1(_00602_),
    .A2(_00612_),
    .B1(_00613_),
    .C1(_00317_),
    .Y(_00614_));
 sky130_fd_sc_hd__inv_2 _07997_ (.A(_06456_),
    .Y(_00615_));
 sky130_fd_sc_hd__a211o_1 _07998_ (.A1(_00317_),
    .A2(_00613_),
    .B1(_00612_),
    .C1(_00602_),
    .X(_00616_));
 sky130_fd_sc_hd__a22o_4 _07999_ (.A1(_03626_),
    .A2(_03928_),
    .B1(_04004_),
    .B2(_03561_),
    .X(_00617_));
 sky130_fd_sc_hd__nand4_2 _08000_ (.A(_00615_),
    .B(_00614_),
    .C(_00616_),
    .D(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__a211oi_1 _08001_ (.A1(_00339_),
    .A2(_00587_),
    .B1(_00586_),
    .C1(_00564_),
    .Y(_00619_));
 sky130_fd_sc_hd__a211o_1 _08002_ (.A1(_00614_),
    .A2(_00618_),
    .B1(_00588_),
    .C1(_00619_),
    .X(_00620_));
 sky130_fd_sc_hd__inv_2 _08003_ (.A(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand3_1 _08004_ (.A(_06508_),
    .B(_06498_),
    .C(_06507_),
    .Y(_00622_));
 sky130_fd_sc_hd__or3_1 _08005_ (.A(_06496_),
    .B(_06490_),
    .C(_06493_),
    .X(_00623_));
 sky130_fd_sc_hd__o21ai_1 _08006_ (.A1(_06496_),
    .A2(_06493_),
    .B1(_06490_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _08007_ (.A(_06488_),
    .B(_05370_),
    .Y(_00625_));
 sky130_fd_sc_hd__a22oi_2 _08008_ (.A1(_06491_),
    .A2(_05434_),
    .B1(_06466_),
    .B2(_06534_),
    .Y(_00626_));
 sky130_fd_sc_hd__and4_1 _08009_ (.A(_02107_),
    .B(_06495_),
    .C(_05434_),
    .D(_06466_),
    .X(_00627_));
 sky130_fd_sc_hd__o21bai_1 _08010_ (.A1(_00625_),
    .A2(_00626_),
    .B1_N(_00627_),
    .Y(_00628_));
 sky130_fd_sc_hd__a21o_1 _08011_ (.A1(_00623_),
    .A2(_00624_),
    .B1(_00628_),
    .X(_00629_));
 sky130_fd_sc_hd__nor2_1 _08012_ (.A(_00531_),
    .B(_00532_),
    .Y(_00630_));
 sky130_fd_sc_hd__xnor2_1 _08013_ (.A(_00529_),
    .B(_00630_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand3_1 _08014_ (.A(_00623_),
    .B(_00628_),
    .C(_00624_),
    .Y(_00632_));
 sky130_fd_sc_hd__a21bo_1 _08015_ (.A1(_00629_),
    .A2(_00631_),
    .B1_N(_00632_),
    .X(_00633_));
 sky130_fd_sc_hd__a21o_1 _08016_ (.A1(_06508_),
    .A2(_06498_),
    .B1(_06507_),
    .X(_00634_));
 sky130_fd_sc_hd__nand3_2 _08017_ (.A(_00622_),
    .B(_00633_),
    .C(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__a21o_1 _08018_ (.A1(_00622_),
    .A2(_00634_),
    .B1(_00633_),
    .X(_00636_));
 sky130_fd_sc_hd__xnor2_1 _08019_ (.A(_00540_),
    .B(_00542_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand3_1 _08020_ (.A(_00635_),
    .B(_00636_),
    .C(_00637_),
    .Y(_00638_));
 sky130_fd_sc_hd__a21oi_2 _08021_ (.A1(_06511_),
    .A2(_06512_),
    .B1(_06532_),
    .Y(_00639_));
 sky130_fd_sc_hd__and3_1 _08022_ (.A(_06511_),
    .B(_06512_),
    .C(_06532_),
    .X(_00640_));
 sky130_fd_sc_hd__a211oi_4 _08023_ (.A1(_00635_),
    .A2(_00638_),
    .B1(_00639_),
    .C1(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hd__o211a_1 _08024_ (.A1(_00640_),
    .A2(_00639_),
    .B1(_00638_),
    .C1(_00635_),
    .X(_00642_));
 sky130_fd_sc_hd__a211o_1 _08025_ (.A1(_00545_),
    .A2(_00560_),
    .B1(_00553_),
    .C1(_00559_),
    .X(_00643_));
 sky130_fd_sc_hd__and4bb_1 _08026_ (.A_N(_00641_),
    .B_N(_00642_),
    .C(_00561_),
    .D(_00643_),
    .X(_00644_));
 sky130_fd_sc_hd__a22o_1 _08027_ (.A1(_06576_),
    .A2(_06577_),
    .B1(_06639_),
    .B2(_06640_),
    .X(_00645_));
 sky130_fd_sc_hd__o211ai_4 _08028_ (.A1(_00641_),
    .A2(_00644_),
    .B1(_00645_),
    .C1(_06641_),
    .Y(_00646_));
 sky130_fd_sc_hd__a211o_1 _08029_ (.A1(_06641_),
    .A2(_00645_),
    .B1(_00644_),
    .C1(_00641_),
    .X(_00647_));
 sky130_fd_sc_hd__a211o_1 _08030_ (.A1(_00579_),
    .A2(_00584_),
    .B1(_00564_),
    .C1(_00585_),
    .X(_00648_));
 sky130_fd_sc_hd__o211ai_2 _08031_ (.A1(_00564_),
    .A2(_00585_),
    .B1(_00579_),
    .C1(_00584_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand4_1 _08032_ (.A(_00646_),
    .B(_00647_),
    .C(_00648_),
    .D(_00649_),
    .Y(_00650_));
 sky130_fd_sc_hd__a22oi_2 _08033_ (.A1(_00026_),
    .A2(_00027_),
    .B1(_00146_),
    .B2(_00147_),
    .Y(_00651_));
 sky130_fd_sc_hd__and4_1 _08034_ (.A(_00026_),
    .B(_00027_),
    .C(_00146_),
    .D(_00147_),
    .X(_00652_));
 sky130_fd_sc_hd__a211o_2 _08035_ (.A1(_00646_),
    .A2(_00650_),
    .B1(_00651_),
    .C1(_00652_),
    .X(_00653_));
 sky130_fd_sc_hd__o211ai_2 _08036_ (.A1(_00652_),
    .A2(_00651_),
    .B1(_00650_),
    .C1(_00646_),
    .Y(_00654_));
 sky130_fd_sc_hd__o211ai_2 _08037_ (.A1(_00588_),
    .A2(_00619_),
    .B1(_00614_),
    .C1(_00618_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand4_2 _08038_ (.A(_00653_),
    .B(_00654_),
    .C(_00620_),
    .D(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__a22oi_2 _08039_ (.A1(_00255_),
    .A2(_00256_),
    .B1(_00368_),
    .B2(_00369_),
    .Y(_00657_));
 sky130_fd_sc_hd__and4_1 _08040_ (.A(_00255_),
    .B(_00256_),
    .C(_00368_),
    .D(_00369_),
    .X(_00658_));
 sky130_fd_sc_hd__a211o_1 _08041_ (.A1(_00653_),
    .A2(_00656_),
    .B1(_00657_),
    .C1(_00658_),
    .X(_00659_));
 sky130_fd_sc_hd__o211ai_1 _08042_ (.A1(_00658_),
    .A2(_00657_),
    .B1(_00656_),
    .C1(_00653_),
    .Y(_00660_));
 sky130_fd_sc_hd__o211a_1 _08043_ (.A1(_00588_),
    .A2(_00621_),
    .B1(_00659_),
    .C1(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__a211oi_2 _08044_ (.A1(_00653_),
    .A2(_00656_),
    .B1(_00657_),
    .C1(_00658_),
    .Y(_00662_));
 sky130_fd_sc_hd__a211o_2 _08045_ (.A1(_00527_),
    .A2(_00528_),
    .B1(_00661_),
    .C1(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__o211ai_4 _08046_ (.A1(_00662_),
    .A2(_00661_),
    .B1(_00528_),
    .C1(_00527_),
    .Y(_00664_));
 sky130_fd_sc_hd__a21boi_2 _08047_ (.A1(_06458_),
    .A2(_00663_),
    .B1_N(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__a31o_1 _08048_ (.A1(_03820_),
    .A2(_03928_),
    .A3(_00516_),
    .B1(_00515_),
    .X(_00666_));
 sky130_fd_sc_hd__or2_1 _08049_ (.A(_00483_),
    .B(_00519_),
    .X(_00667_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_00483_),
    .B(_00519_),
    .Y(_00668_));
 sky130_fd_sc_hd__a21bo_2 _08051_ (.A1(_00482_),
    .A2(_00667_),
    .B1_N(_00668_),
    .X(_00669_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(_00499_),
    .B(_00500_),
    .Y(_00670_));
 sky130_fd_sc_hd__or2_1 _08053_ (.A(_00499_),
    .B(_00500_),
    .X(_00671_));
 sky130_fd_sc_hd__a21boi_4 _08054_ (.A1(_00670_),
    .A2(_00518_),
    .B1_N(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__o21bai_2 _08055_ (.A1(_00441_),
    .A2(_00475_),
    .B1_N(_00474_),
    .Y(_00673_));
 sky130_fd_sc_hd__or3_1 _08056_ (.A(_00509_),
    .B(_00510_),
    .C(_00512_),
    .X(_00674_));
 sky130_fd_sc_hd__or2b_1 _08057_ (.A(_00505_),
    .B_N(_00513_),
    .X(_00675_));
 sky130_fd_sc_hd__buf_2 _08058_ (.A(_03593_),
    .X(_00676_));
 sky130_fd_sc_hd__a22oi_1 _08059_ (.A1(_00676_),
    .A2(_04176_),
    .B1(_04240_),
    .B2(_00506_),
    .Y(_00677_));
 sky130_fd_sc_hd__clkbuf_2 _08060_ (.A(net57),
    .X(_00678_));
 sky130_fd_sc_hd__and4_1 _08061_ (.A(_03539_),
    .B(_00678_),
    .C(_00287_),
    .D(_00267_),
    .X(_00679_));
 sky130_fd_sc_hd__nor2_1 _08062_ (.A(_00677_),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _08063_ (.A(_06439_),
    .B(_00303_),
    .Y(_00681_));
 sky130_fd_sc_hd__xnor2_1 _08064_ (.A(_00680_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_1 _08065_ (.A(_00508_),
    .B(_00509_),
    .Y(_00683_));
 sky130_fd_sc_hd__xnor2_1 _08066_ (.A(_00682_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2_1 _08067_ (.A(_06429_),
    .B(_04057_),
    .Y(_00685_));
 sky130_fd_sc_hd__xor2_1 _08068_ (.A(_00684_),
    .B(_00685_),
    .X(_00686_));
 sky130_fd_sc_hd__a21oi_1 _08069_ (.A1(_00674_),
    .A2(_00675_),
    .B1(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__and3_1 _08070_ (.A(_00674_),
    .B(_00675_),
    .C(_00686_),
    .X(_00688_));
 sky130_fd_sc_hd__nor2_2 _08071_ (.A(_00687_),
    .B(_00688_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_00502_),
    .B(_03993_),
    .Y(_00690_));
 sky130_fd_sc_hd__xnor2_4 _08073_ (.A(_00689_),
    .B(_00690_),
    .Y(_00691_));
 sky130_fd_sc_hd__a21o_1 _08074_ (.A1(_00460_),
    .A2(_00469_),
    .B1(_00468_),
    .X(_00692_));
 sky130_fd_sc_hd__a32o_1 _08075_ (.A1(_00270_),
    .A2(_00093_),
    .A3(_00457_),
    .B1(_00230_),
    .B2(_00036_),
    .X(_00693_));
 sky130_fd_sc_hd__a22o_1 _08076_ (.A1(_03432_),
    .A2(_04358_),
    .B1(_00083_),
    .B2(_00278_),
    .X(_00694_));
 sky130_fd_sc_hd__nand4_2 _08077_ (.A(_03378_),
    .B(_00279_),
    .C(_04358_),
    .D(_00083_),
    .Y(_00695_));
 sky130_fd_sc_hd__a22o_1 _08078_ (.A1(_00292_),
    .A2(_00259_),
    .B1(_00694_),
    .B2(_00695_),
    .X(_00696_));
 sky130_fd_sc_hd__nand4_2 _08079_ (.A(_00283_),
    .B(_00259_),
    .C(_00694_),
    .D(_00695_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3_2 _08080_ (.A(_00693_),
    .B(_00696_),
    .C(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__a21o_1 _08081_ (.A1(_00696_),
    .A2(_00697_),
    .B1(_00693_),
    .X(_00699_));
 sky130_fd_sc_hd__nand2_1 _08082_ (.A(_00488_),
    .B(_00490_),
    .Y(_00700_));
 sky130_fd_sc_hd__a21o_1 _08083_ (.A1(_00698_),
    .A2(_00699_),
    .B1(_00700_),
    .X(_00701_));
 sky130_fd_sc_hd__nand3_2 _08084_ (.A(_00700_),
    .B(_00698_),
    .C(_00699_),
    .Y(_00702_));
 sky130_fd_sc_hd__and3_1 _08085_ (.A(_00692_),
    .B(_00701_),
    .C(_00702_),
    .X(_00703_));
 sky130_fd_sc_hd__a21oi_1 _08086_ (.A1(_00701_),
    .A2(_00702_),
    .B1(_00692_),
    .Y(_00704_));
 sky130_fd_sc_hd__a211oi_1 _08087_ (.A1(_00491_),
    .A2(_00493_),
    .B1(_00703_),
    .C1(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__o211a_1 _08088_ (.A1(_00703_),
    .A2(_00704_),
    .B1(_00491_),
    .C1(_00493_),
    .X(_00706_));
 sky130_fd_sc_hd__or2_2 _08089_ (.A(_00705_),
    .B(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__nor2_2 _08090_ (.A(_00495_),
    .B(_00497_),
    .Y(_00708_));
 sky130_fd_sc_hd__xnor2_1 _08091_ (.A(_00707_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__xnor2_1 _08092_ (.A(_00691_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__xnor2_2 _08093_ (.A(_00673_),
    .B(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__xor2_2 _08094_ (.A(_00672_),
    .B(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__nor2_2 _08095_ (.A(_00455_),
    .B(_00472_),
    .Y(_00713_));
 sky130_fd_sc_hd__o21bai_1 _08096_ (.A1(_00422_),
    .A2(_00424_),
    .B1_N(_00425_),
    .Y(_00714_));
 sky130_fd_sc_hd__a22o_1 _08097_ (.A1(_00062_),
    .A2(_06591_),
    .B1(_06584_),
    .B2(_00049_),
    .X(_00715_));
 sky130_fd_sc_hd__nand4_1 _08098_ (.A(_00217_),
    .B(_00216_),
    .C(_06591_),
    .D(_05036_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand4_1 _08099_ (.A(_00221_),
    .B(_04918_),
    .C(_00715_),
    .D(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__a22o_1 _08100_ (.A1(_00444_),
    .A2(_00550_),
    .B1(_00715_),
    .B2(_00716_),
    .X(_00718_));
 sky130_fd_sc_hd__nand3_1 _08101_ (.A(_00714_),
    .B(_00717_),
    .C(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__a21o_1 _08102_ (.A1(_00717_),
    .A2(_00718_),
    .B1(_00714_),
    .X(_00720_));
 sky130_fd_sc_hd__nand2_1 _08103_ (.A(_00447_),
    .B(_00449_),
    .Y(_00721_));
 sky130_fd_sc_hd__a21o_1 _08104_ (.A1(_00719_),
    .A2(_00720_),
    .B1(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__nand3_1 _08105_ (.A(_00721_),
    .B(_00719_),
    .C(_00720_),
    .Y(_00723_));
 sky130_fd_sc_hd__a21bo_1 _08106_ (.A1(_00442_),
    .A2(_00451_),
    .B1_N(_00450_),
    .X(_00724_));
 sky130_fd_sc_hd__and3_1 _08107_ (.A(_00722_),
    .B(_00723_),
    .C(_00724_),
    .X(_00725_));
 sky130_fd_sc_hd__a21oi_1 _08108_ (.A1(_00722_),
    .A2(_00723_),
    .B1(_00724_),
    .Y(_00726_));
 sky130_fd_sc_hd__buf_4 _08109_ (.A(_00231_),
    .X(_00727_));
 sky130_fd_sc_hd__buf_4 _08110_ (.A(_00299_),
    .X(_00728_));
 sky130_fd_sc_hd__a22oi_1 _08111_ (.A1(_00727_),
    .A2(_00036_),
    .B1(_00059_),
    .B2(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__and4_1 _08112_ (.A(_03228_),
    .B(_03282_),
    .C(_04585_),
    .D(_04649_),
    .X(_00730_));
 sky130_fd_sc_hd__nor2_1 _08113_ (.A(_00729_),
    .B(_00730_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _08114_ (.A(_00077_),
    .B(_04531_),
    .Y(_00732_));
 sky130_fd_sc_hd__xnor2_1 _08115_ (.A(_00731_),
    .B(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__a22oi_4 _08116_ (.A1(_03099_),
    .A2(_04778_),
    .B1(_06603_),
    .B2(_03056_),
    .Y(_00734_));
 sky130_fd_sc_hd__and4_1 _08117_ (.A(_00237_),
    .B(_00462_),
    .C(_04778_),
    .D(_04832_),
    .X(_00735_));
 sky130_fd_sc_hd__nand2_1 _08118_ (.A(_00088_),
    .B(_00040_),
    .Y(_00736_));
 sky130_fd_sc_hd__or3_1 _08119_ (.A(_00734_),
    .B(_00735_),
    .C(_00736_),
    .X(_00737_));
 sky130_fd_sc_hd__o21ai_1 _08120_ (.A1(_00734_),
    .A2(_00735_),
    .B1(_00736_),
    .Y(_00738_));
 sky130_fd_sc_hd__o21bai_2 _08121_ (.A1(_00461_),
    .A2(_00463_),
    .B1_N(_00464_),
    .Y(_00739_));
 sky130_fd_sc_hd__and3_1 _08122_ (.A(_00737_),
    .B(_00738_),
    .C(_00739_),
    .X(_00740_));
 sky130_fd_sc_hd__a21o_1 _08123_ (.A1(_00737_),
    .A2(_00738_),
    .B1(_00739_),
    .X(_00741_));
 sky130_fd_sc_hd__or2b_1 _08124_ (.A(_00740_),
    .B_N(_00741_),
    .X(_00742_));
 sky130_fd_sc_hd__xnor2_1 _08125_ (.A(_00733_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__o21ba_1 _08126_ (.A1(_00725_),
    .A2(_00726_),
    .B1_N(_00743_),
    .X(_00744_));
 sky130_fd_sc_hd__nor3b_1 _08127_ (.A(_00725_),
    .B(_00726_),
    .C_N(_00743_),
    .Y(_00745_));
 sky130_fd_sc_hd__a211o_1 _08128_ (.A1(_00430_),
    .A2(_00433_),
    .B1(_00744_),
    .C1(_00745_),
    .X(_00746_));
 sky130_fd_sc_hd__o211ai_1 _08129_ (.A1(_00744_),
    .A2(_00745_),
    .B1(_00430_),
    .C1(_00433_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(_00746_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__xor2_2 _08131_ (.A(_00713_),
    .B(_00748_),
    .X(_00749_));
 sky130_fd_sc_hd__a21o_1 _08132_ (.A1(_00394_),
    .A2(_00403_),
    .B1(_00402_),
    .X(_00750_));
 sky130_fd_sc_hd__a22oi_1 _08133_ (.A1(_06601_),
    .A2(_05187_),
    .B1(_06568_),
    .B2(_06606_),
    .Y(_00751_));
 sky130_fd_sc_hd__and4_1 _08134_ (.A(_02754_),
    .B(_02797_),
    .C(_05187_),
    .D(_06518_),
    .X(_00752_));
 sky130_fd_sc_hd__nor2_1 _08135_ (.A(_00751_),
    .B(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _08136_ (.A(_02840_),
    .B(_00423_),
    .Y(_00754_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(_00753_),
    .B(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__a22oi_2 _08138_ (.A1(_06622_),
    .A2(_05370_),
    .B1(_06489_),
    .B2(_00414_),
    .Y(_00756_));
 sky130_fd_sc_hd__and4_1 _08139_ (.A(_06578_),
    .B(_06579_),
    .C(_05370_),
    .D(_05434_),
    .X(_00757_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(net122),
    .B(_06562_),
    .Y(_00758_));
 sky130_fd_sc_hd__or3_1 _08141_ (.A(_00756_),
    .B(_00757_),
    .C(_00758_),
    .X(_00759_));
 sky130_fd_sc_hd__o21ai_1 _08142_ (.A1(_00756_),
    .A2(_00757_),
    .B1(_00758_),
    .Y(_00760_));
 sky130_fd_sc_hd__o21bai_1 _08143_ (.A1(_00411_),
    .A2(_00413_),
    .B1_N(_00415_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand3_2 _08144_ (.A(_00759_),
    .B(_00760_),
    .C(_00761_),
    .Y(_00762_));
 sky130_fd_sc_hd__a21o_1 _08145_ (.A1(_00759_),
    .A2(_00760_),
    .B1(_00761_),
    .X(_00763_));
 sky130_fd_sc_hd__nand3_1 _08146_ (.A(_00755_),
    .B(_00762_),
    .C(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__a21o_1 _08147_ (.A1(_00762_),
    .A2(_00763_),
    .B1(_00755_),
    .X(_00765_));
 sky130_fd_sc_hd__and3_1 _08148_ (.A(_00750_),
    .B(_00764_),
    .C(_00765_),
    .X(_00766_));
 sky130_fd_sc_hd__a21oi_1 _08149_ (.A1(_00764_),
    .A2(_00765_),
    .B1(_00750_),
    .Y(_00767_));
 sky130_fd_sc_hd__a211o_1 _08150_ (.A1(_00419_),
    .A2(_00428_),
    .B1(_00766_),
    .C1(_00767_),
    .X(_00768_));
 sky130_fd_sc_hd__o211ai_1 _08151_ (.A1(_00766_),
    .A2(_00767_),
    .B1(_00419_),
    .C1(_00428_),
    .Y(_00769_));
 sky130_fd_sc_hd__and2_1 _08152_ (.A(_00768_),
    .B(_00769_),
    .X(_00770_));
 sky130_fd_sc_hd__nand2_1 _08153_ (.A(_00399_),
    .B(_00400_),
    .Y(_00771_));
 sky130_fd_sc_hd__o21bai_1 _08154_ (.A1(_00383_),
    .A2(_00386_),
    .B1_N(_00384_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_06663_),
    .B(_00398_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand4_1 _08156_ (.A(_06565_),
    .B(_06516_),
    .C(_05563_),
    .D(_05638_),
    .Y(_00774_));
 sky130_fd_sc_hd__a22o_1 _08157_ (.A1(_06516_),
    .A2(_06461_),
    .B1(_05638_),
    .B2(_06520_),
    .X(_00775_));
 sky130_fd_sc_hd__nand3b_1 _08158_ (.A_N(_00773_),
    .B(_00774_),
    .C(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__a21bo_1 _08159_ (.A1(_00775_),
    .A2(_00774_),
    .B1_N(_00773_),
    .X(_00777_));
 sky130_fd_sc_hd__and3_1 _08160_ (.A(_00772_),
    .B(_00776_),
    .C(_00777_),
    .X(_00778_));
 sky130_fd_sc_hd__a21o_1 _08161_ (.A1(_00776_),
    .A2(_00777_),
    .B1(_00772_),
    .X(_00779_));
 sky130_fd_sc_hd__and2b_1 _08162_ (.A_N(_00778_),
    .B(_00779_),
    .X(_00780_));
 sky130_fd_sc_hd__xnor2_2 _08163_ (.A(_00771_),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(_02377_),
    .B(_05702_),
    .Y(_00782_));
 sky130_fd_sc_hd__clkbuf_4 _08165_ (.A(net128),
    .X(_00783_));
 sky130_fd_sc_hd__a22oi_1 _08166_ (.A1(_00162_),
    .A2(_05756_),
    .B1(_00783_),
    .B2(_00164_),
    .Y(_00784_));
 sky130_fd_sc_hd__buf_2 _08167_ (.A(net128),
    .X(_00785_));
 sky130_fd_sc_hd__and4_1 _08168_ (.A(_06501_),
    .B(_06500_),
    .C(_05756_),
    .D(_00785_),
    .X(_00786_));
 sky130_fd_sc_hd__nor2_1 _08169_ (.A(_00784_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__xnor2_2 _08170_ (.A(_00782_),
    .B(_00787_),
    .Y(_00788_));
 sky130_fd_sc_hd__clkbuf_4 _08171_ (.A(net29),
    .X(_00789_));
 sky130_fd_sc_hd__a22oi_1 _08172_ (.A1(_02248_),
    .A2(_00153_),
    .B1(_00789_),
    .B2(_02205_),
    .Y(_00790_));
 sky130_fd_sc_hd__and4_1 _08173_ (.A(_06463_),
    .B(net111),
    .C(net28),
    .D(net29),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _08174_ (.A(_00790_),
    .B(_00791_),
    .X(_00792_));
 sky130_fd_sc_hd__a21bo_1 _08175_ (.A1(_00375_),
    .A2(_00376_),
    .B1_N(_00374_),
    .X(_00793_));
 sky130_fd_sc_hd__xnor2_2 _08176_ (.A(_00792_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__xnor2_2 _08177_ (.A(_00788_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__a21bo_1 _08178_ (.A1(_00381_),
    .A2(_00388_),
    .B1_N(_00380_),
    .X(_00796_));
 sky130_fd_sc_hd__xor2_2 _08179_ (.A(_00795_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__xnor2_2 _08180_ (.A(_00781_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__a21bo_1 _08181_ (.A1(_00393_),
    .A2(_00405_),
    .B1_N(_00392_),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_1 _08182_ (.A(_00798_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__xnor2_1 _08183_ (.A(_00770_),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__a21bo_1 _08184_ (.A1(_00409_),
    .A2(_00435_),
    .B1_N(_00408_),
    .X(_00802_));
 sky130_fd_sc_hd__xnor2_1 _08185_ (.A(_00801_),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__xor2_2 _08186_ (.A(_00749_),
    .B(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__a21boi_1 _08187_ (.A1(_00439_),
    .A2(_00477_),
    .B1_N(_00438_),
    .Y(_00805_));
 sky130_fd_sc_hd__xnor2_2 _08188_ (.A(_00804_),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__xnor2_2 _08189_ (.A(_00712_),
    .B(_00806_),
    .Y(_00807_));
 sky130_fd_sc_hd__a21boi_2 _08190_ (.A1(_00481_),
    .A2(_00521_),
    .B1_N(_00480_),
    .Y(_00808_));
 sky130_fd_sc_hd__xnor2_2 _08191_ (.A(_00807_),
    .B(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hd__xor2_4 _08192_ (.A(_00669_),
    .B(_00809_),
    .X(_00810_));
 sky130_fd_sc_hd__a21boi_4 _08193_ (.A1(_00525_),
    .A2(_00526_),
    .B1_N(_00524_),
    .Y(_00811_));
 sky130_fd_sc_hd__xor2_2 _08194_ (.A(_00810_),
    .B(_00811_),
    .X(_00812_));
 sky130_fd_sc_hd__xor2_1 _08195_ (.A(_00666_),
    .B(_00812_),
    .X(_00813_));
 sky130_fd_sc_hd__and2b_1 _08196_ (.A_N(_00665_),
    .B(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__or2b_1 _08197_ (.A(_00813_),
    .B_N(_00665_),
    .X(_00815_));
 sky130_fd_sc_hd__or2b_1 _08198_ (.A(_00814_),
    .B_N(_00815_),
    .X(_00816_));
 sky130_fd_sc_hd__nand3_1 _08199_ (.A(_06458_),
    .B(_00664_),
    .C(_00663_),
    .Y(_00817_));
 sky130_fd_sc_hd__a21o_1 _08200_ (.A1(_00664_),
    .A2(_00663_),
    .B1(_06458_),
    .X(_00818_));
 sky130_fd_sc_hd__nand3_1 _08201_ (.A(_00632_),
    .B(_00629_),
    .C(_00631_),
    .Y(_00819_));
 sky130_fd_sc_hd__a22oi_2 _08202_ (.A1(_00162_),
    .A2(_06518_),
    .B1(_00412_),
    .B2(_00164_),
    .Y(_00820_));
 sky130_fd_sc_hd__and4_1 _08203_ (.A(_06501_),
    .B(_06548_),
    .C(_05241_),
    .D(_06562_),
    .X(_00821_));
 sky130_fd_sc_hd__nor2_1 _08204_ (.A(_00820_),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(_06475_),
    .B(_06525_),
    .Y(_00823_));
 sky130_fd_sc_hd__xnor2_1 _08206_ (.A(_00822_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__or3_1 _08207_ (.A(_00627_),
    .B(_00625_),
    .C(_00626_),
    .X(_00825_));
 sky130_fd_sc_hd__o21ai_1 _08208_ (.A1(_00627_),
    .A2(_00626_),
    .B1(_00625_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(_06460_),
    .B(_05305_),
    .Y(_00827_));
 sky130_fd_sc_hd__a22oi_2 _08210_ (.A1(_06463_),
    .A2(net19),
    .B1(_05434_),
    .B2(_02107_),
    .Y(_00828_));
 sky130_fd_sc_hd__and4_1 _08211_ (.A(_06469_),
    .B(_02194_),
    .C(net19),
    .D(net20),
    .X(_00829_));
 sky130_fd_sc_hd__o21bai_1 _08212_ (.A1(_00827_),
    .A2(_00828_),
    .B1_N(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__a21o_1 _08213_ (.A1(_00825_),
    .A2(_00826_),
    .B1(_00830_),
    .X(_00831_));
 sky130_fd_sc_hd__nand3_1 _08214_ (.A(_00825_),
    .B(_00830_),
    .C(_00826_),
    .Y(_00832_));
 sky130_fd_sc_hd__a21bo_1 _08215_ (.A1(_00824_),
    .A2(_00831_),
    .B1_N(_00832_),
    .X(_00833_));
 sky130_fd_sc_hd__a21o_1 _08216_ (.A1(_00632_),
    .A2(_00629_),
    .B1(_00631_),
    .X(_00834_));
 sky130_fd_sc_hd__nand3_4 _08217_ (.A(_00819_),
    .B(_00833_),
    .C(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__o21ba_1 _08218_ (.A1(_00820_),
    .A2(_00823_),
    .B1_N(_00821_),
    .X(_00836_));
 sky130_fd_sc_hd__o2bb2a_1 _08219_ (.A1_N(_02528_),
    .A2_N(_05036_),
    .B1(_00537_),
    .B2(_00538_),
    .X(_00837_));
 sky130_fd_sc_hd__nor2_1 _08220_ (.A(_00539_),
    .B(_00837_),
    .Y(_00838_));
 sky130_fd_sc_hd__xnor2_1 _08221_ (.A(_00836_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand2_1 _08222_ (.A(_06560_),
    .B(_04972_),
    .Y(_00840_));
 sky130_fd_sc_hd__a22oi_2 _08223_ (.A1(_02485_),
    .A2(_06584_),
    .B1(_05112_),
    .B2(_06565_),
    .Y(_00841_));
 sky130_fd_sc_hd__and4_1 _08224_ (.A(_02420_),
    .B(_06513_),
    .C(_05025_),
    .D(_05101_),
    .X(_00842_));
 sky130_fd_sc_hd__o21ba_1 _08225_ (.A1(_00840_),
    .A2(_00841_),
    .B1_N(_00842_),
    .X(_00843_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_00839_),
    .B(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__a21o_1 _08227_ (.A1(_00819_),
    .A2(_00834_),
    .B1(_00833_),
    .X(_00845_));
 sky130_fd_sc_hd__nand3_2 _08228_ (.A(_00835_),
    .B(_00844_),
    .C(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__a21oi_2 _08229_ (.A1(_00635_),
    .A2(_00636_),
    .B1(_00637_),
    .Y(_00847_));
 sky130_fd_sc_hd__and3_1 _08230_ (.A(_00635_),
    .B(_00636_),
    .C(_00637_),
    .X(_00848_));
 sky130_fd_sc_hd__a211oi_4 _08231_ (.A1(_00835_),
    .A2(_00846_),
    .B1(_00847_),
    .C1(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__o2bb2a_1 _08232_ (.A1_N(_06620_),
    .A2_N(_00445_),
    .B1(_00546_),
    .B2(_00547_),
    .X(_00850_));
 sky130_fd_sc_hd__nor2_1 _08233_ (.A(_00548_),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__and4_1 _08234_ (.A(_06578_),
    .B(_02647_),
    .C(_06602_),
    .D(_06604_),
    .X(_00852_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(net122),
    .B(_04778_),
    .Y(_00853_));
 sky130_fd_sc_hd__a22oi_2 _08236_ (.A1(_06622_),
    .A2(_04832_),
    .B1(_04896_),
    .B2(_00414_),
    .Y(_00854_));
 sky130_fd_sc_hd__or3_1 _08237_ (.A(_00852_),
    .B(_00853_),
    .C(_00854_),
    .X(_00855_));
 sky130_fd_sc_hd__or2b_1 _08238_ (.A(_00852_),
    .B_N(_00855_),
    .X(_00856_));
 sky130_fd_sc_hd__and2_1 _08239_ (.A(_00851_),
    .B(_00856_),
    .X(_00857_));
 sky130_fd_sc_hd__xor2_1 _08240_ (.A(_00851_),
    .B(_00856_),
    .X(_00858_));
 sky130_fd_sc_hd__nand2_1 _08241_ (.A(_02851_),
    .B(_04660_),
    .Y(_00859_));
 sky130_fd_sc_hd__a21boi_2 _08242_ (.A1(_00555_),
    .A2(_00566_),
    .B1_N(_00565_),
    .Y(_00860_));
 sky130_fd_sc_hd__xnor2_2 _08243_ (.A(_00859_),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__and2_1 _08244_ (.A(_00858_),
    .B(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__or3_1 _08245_ (.A(_00539_),
    .B(_00836_),
    .C(_00837_),
    .X(_00863_));
 sky130_fd_sc_hd__or2b_1 _08246_ (.A(_00843_),
    .B_N(_00839_),
    .X(_00864_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(_00554_),
    .B(_00558_),
    .Y(_00865_));
 sky130_fd_sc_hd__a21o_2 _08248_ (.A1(_00863_),
    .A2(_00864_),
    .B1(_00865_),
    .X(_00866_));
 sky130_fd_sc_hd__nand3_1 _08249_ (.A(_00863_),
    .B(_00864_),
    .C(_00865_),
    .Y(_00867_));
 sky130_fd_sc_hd__o211ai_4 _08250_ (.A1(_00857_),
    .A2(_00862_),
    .B1(_00866_),
    .C1(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__a211o_1 _08251_ (.A1(_00866_),
    .A2(_00867_),
    .B1(_00857_),
    .C1(_00862_),
    .X(_00869_));
 sky130_fd_sc_hd__o211ai_1 _08252_ (.A1(_00848_),
    .A2(_00847_),
    .B1(_00846_),
    .C1(_00835_),
    .Y(_00870_));
 sky130_fd_sc_hd__and4b_2 _08253_ (.A_N(_00849_),
    .B(_00868_),
    .C(_00869_),
    .D(_00870_),
    .X(_00871_));
 sky130_fd_sc_hd__a2bb2o_1 _08254_ (.A1_N(_00641_),
    .A2_N(_00642_),
    .B1(_00561_),
    .B2(_00643_),
    .X(_00872_));
 sky130_fd_sc_hd__or4bb_2 _08255_ (.A(_00641_),
    .B(_00642_),
    .C_N(_00561_),
    .D_N(_00643_),
    .X(_00873_));
 sky130_fd_sc_hd__o211ai_4 _08256_ (.A1(_00849_),
    .A2(_00871_),
    .B1(_00872_),
    .C1(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__and2_1 _08257_ (.A(net121),
    .B(_04585_),
    .X(_00875_));
 sky130_fd_sc_hd__a22o_1 _08258_ (.A1(_00011_),
    .A2(_00048_),
    .B1(_00040_),
    .B2(_00012_),
    .X(_00876_));
 sky130_fd_sc_hd__buf_4 _08259_ (.A(_06598_),
    .X(_00877_));
 sky130_fd_sc_hd__buf_4 _08260_ (.A(_06599_),
    .X(_00878_));
 sky130_fd_sc_hd__nand4_2 _08261_ (.A(_00877_),
    .B(_00878_),
    .C(_04649_),
    .D(_04714_),
    .Y(_00879_));
 sky130_fd_sc_hd__a21bo_1 _08262_ (.A1(_00875_),
    .A2(_00876_),
    .B1_N(_00879_),
    .X(_00880_));
 sky130_fd_sc_hd__o21ai_1 _08263_ (.A1(_00571_),
    .A2(_00573_),
    .B1(_00572_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand3_1 _08264_ (.A(_00574_),
    .B(_00880_),
    .C(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__and4_1 _08265_ (.A(_02894_),
    .B(_02948_),
    .C(_00083_),
    .D(_00098_),
    .X(_00883_));
 sky130_fd_sc_hd__nand2_1 _08266_ (.A(net119),
    .B(_00090_),
    .Y(_00884_));
 sky130_fd_sc_hd__a22oi_1 _08267_ (.A1(_00062_),
    .A2(_04445_),
    .B1(_00085_),
    .B2(_00063_),
    .Y(_00885_));
 sky130_fd_sc_hd__or3_1 _08268_ (.A(_00883_),
    .B(_00884_),
    .C(_00885_),
    .X(_00886_));
 sky130_fd_sc_hd__or2b_1 _08269_ (.A(_00883_),
    .B_N(_00886_),
    .X(_00887_));
 sky130_fd_sc_hd__a21o_1 _08270_ (.A1(_00574_),
    .A2(_00881_),
    .B1(_00880_),
    .X(_00888_));
 sky130_fd_sc_hd__nand3_1 _08271_ (.A(_00882_),
    .B(_00887_),
    .C(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__xnor2_1 _08272_ (.A(_00575_),
    .B(_00576_),
    .Y(_00890_));
 sky130_fd_sc_hd__a21o_1 _08273_ (.A1(_00882_),
    .A2(_00889_),
    .B1(_00890_),
    .X(_00891_));
 sky130_fd_sc_hd__a21oi_1 _08274_ (.A1(_00882_),
    .A2(_00889_),
    .B1(_00890_),
    .Y(_00892_));
 sky130_fd_sc_hd__and3_1 _08275_ (.A(_00890_),
    .B(_00882_),
    .C(_00889_),
    .X(_00893_));
 sky130_fd_sc_hd__and3_1 _08276_ (.A(_00599_),
    .B(_00590_),
    .C(_00598_),
    .X(_00894_));
 sky130_fd_sc_hd__a21oi_1 _08277_ (.A1(_00599_),
    .A2(_00598_),
    .B1(_00590_),
    .Y(_00895_));
 sky130_fd_sc_hd__or2_2 _08278_ (.A(_00894_),
    .B(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__or3_1 _08279_ (.A(_00892_),
    .B(_00893_),
    .C(_00896_),
    .X(_00897_));
 sky130_fd_sc_hd__o21a_1 _08280_ (.A1(_00580_),
    .A2(_00581_),
    .B1(_00583_),
    .X(_00898_));
 sky130_fd_sc_hd__nor3_2 _08281_ (.A(_00580_),
    .B(_00581_),
    .C(_00583_),
    .Y(_00899_));
 sky130_fd_sc_hd__a211oi_4 _08282_ (.A1(_00866_),
    .A2(_00868_),
    .B1(_00898_),
    .C1(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__o211a_1 _08283_ (.A1(_00899_),
    .A2(_00898_),
    .B1(_00868_),
    .C1(_00866_),
    .X(_00901_));
 sky130_fd_sc_hd__a211o_1 _08284_ (.A1(_00891_),
    .A2(_00897_),
    .B1(_00900_),
    .C1(_00901_),
    .X(_00902_));
 sky130_fd_sc_hd__o211ai_2 _08285_ (.A1(_00900_),
    .A2(_00901_),
    .B1(_00891_),
    .C1(_00897_),
    .Y(_00903_));
 sky130_fd_sc_hd__a211o_1 _08286_ (.A1(_00873_),
    .A2(_00872_),
    .B1(_00871_),
    .C1(_00849_),
    .X(_00904_));
 sky130_fd_sc_hd__nand4_1 _08287_ (.A(_00874_),
    .B(_00902_),
    .C(_00903_),
    .D(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__a22oi_2 _08288_ (.A1(_00646_),
    .A2(_00647_),
    .B1(_00648_),
    .B2(_00649_),
    .Y(_00906_));
 sky130_fd_sc_hd__and4_1 _08289_ (.A(_00646_),
    .B(_00647_),
    .C(_00648_),
    .D(_00649_),
    .X(_00907_));
 sky130_fd_sc_hd__a211o_1 _08290_ (.A1(_00874_),
    .A2(_00905_),
    .B1(_00906_),
    .C1(_00907_),
    .X(_00908_));
 sky130_fd_sc_hd__xnor2_1 _08291_ (.A(_00610_),
    .B(_00611_),
    .Y(_00909_));
 sky130_fd_sc_hd__a22oi_1 _08292_ (.A1(_03454_),
    .A2(_03884_),
    .B1(_03982_),
    .B2(_03389_),
    .Y(_00910_));
 sky130_fd_sc_hd__or2_1 _08293_ (.A(_00608_),
    .B(_00910_),
    .X(_00911_));
 sky130_fd_sc_hd__a22o_1 _08294_ (.A1(_03293_),
    .A2(_04046_),
    .B1(_04122_),
    .B2(_03239_),
    .X(_00912_));
 sky130_fd_sc_hd__and4_1 _08295_ (.A(_00728_),
    .B(_00727_),
    .C(_04046_),
    .D(_00303_),
    .X(_00913_));
 sky130_fd_sc_hd__a31o_1 _08296_ (.A1(_03346_),
    .A2(_03982_),
    .A3(_00912_),
    .B1(_00913_),
    .X(_00914_));
 sky130_fd_sc_hd__and2b_2 _08297_ (.A_N(_00911_),
    .B(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__nand2_1 _08298_ (.A(_03335_),
    .B(_04057_),
    .Y(_00916_));
 sky130_fd_sc_hd__and2b_1 _08299_ (.A_N(_00605_),
    .B(_00604_),
    .X(_00917_));
 sky130_fd_sc_hd__xnor2_2 _08300_ (.A(_00916_),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__o21ai_2 _08301_ (.A1(_00593_),
    .A2(_00595_),
    .B1(_00594_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _08302_ (.A(_00262_),
    .B(_00272_),
    .Y(_00920_));
 sky130_fd_sc_hd__buf_6 _08303_ (.A(_00237_),
    .X(_00921_));
 sky130_fd_sc_hd__a22oi_4 _08304_ (.A1(_03110_),
    .A2(_00301_),
    .B1(_00259_),
    .B2(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__and4_1 _08305_ (.A(_00133_),
    .B(_00132_),
    .C(_04240_),
    .D(_04305_),
    .X(_00923_));
 sky130_fd_sc_hd__o21bai_1 _08306_ (.A1(_00920_),
    .A2(_00922_),
    .B1_N(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__a21o_1 _08307_ (.A1(_00596_),
    .A2(_00919_),
    .B1(_00924_),
    .X(_00925_));
 sky130_fd_sc_hd__and3_1 _08308_ (.A(_00596_),
    .B(_00919_),
    .C(_00924_),
    .X(_00926_));
 sky130_fd_sc_hd__a21oi_1 _08309_ (.A1(_00918_),
    .A2(_00925_),
    .B1(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__or2b_1 _08310_ (.A(_00609_),
    .B_N(_00607_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_2 _08311_ (.A(_00928_),
    .B(_00608_),
    .Y(_00929_));
 sky130_fd_sc_hd__xnor2_1 _08312_ (.A(_00927_),
    .B(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__and2b_1 _08313_ (.A_N(_00927_),
    .B(_00929_),
    .X(_00931_));
 sky130_fd_sc_hd__a21oi_1 _08314_ (.A1(_00915_),
    .A2(_00930_),
    .B1(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__or2_1 _08315_ (.A(_00909_),
    .B(_00932_),
    .X(_00933_));
 sky130_fd_sc_hd__nand2_2 _08316_ (.A(_03561_),
    .B(_03928_),
    .Y(_00934_));
 sky130_fd_sc_hd__xnor2_1 _08317_ (.A(_00909_),
    .B(_00932_),
    .Y(_00935_));
 sky130_fd_sc_hd__or2_1 _08318_ (.A(_00934_),
    .B(_00935_),
    .X(_00936_));
 sky130_fd_sc_hd__a211oi_1 _08319_ (.A1(_00891_),
    .A2(_00897_),
    .B1(_00900_),
    .C1(_00901_),
    .Y(_00937_));
 sky130_fd_sc_hd__a22o_1 _08320_ (.A1(_00614_),
    .A2(_00616_),
    .B1(_00617_),
    .B2(_00615_),
    .X(_00938_));
 sky130_fd_sc_hd__o211a_1 _08321_ (.A1(_00900_),
    .A2(_00937_),
    .B1(_00938_),
    .C1(_00618_),
    .X(_00939_));
 sky130_fd_sc_hd__a211oi_1 _08322_ (.A1(_00618_),
    .A2(_00938_),
    .B1(_00937_),
    .C1(_00900_),
    .Y(_00940_));
 sky130_fd_sc_hd__a211o_1 _08323_ (.A1(_00933_),
    .A2(_00936_),
    .B1(_00939_),
    .C1(_00940_),
    .X(_00941_));
 sky130_fd_sc_hd__o211ai_2 _08324_ (.A1(_00939_),
    .A2(_00940_),
    .B1(_00933_),
    .C1(_00936_),
    .Y(_00942_));
 sky130_fd_sc_hd__o211ai_2 _08325_ (.A1(_00907_),
    .A2(_00906_),
    .B1(_00905_),
    .C1(_00874_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand4_1 _08326_ (.A(_00908_),
    .B(_00941_),
    .C(_00942_),
    .D(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__a22oi_2 _08327_ (.A1(_00653_),
    .A2(_00654_),
    .B1(_00620_),
    .B2(_00655_),
    .Y(_00945_));
 sky130_fd_sc_hd__and4_1 _08328_ (.A(_00653_),
    .B(_00654_),
    .C(_00620_),
    .D(_00655_),
    .X(_00946_));
 sky130_fd_sc_hd__a211oi_1 _08329_ (.A1(_00908_),
    .A2(_00944_),
    .B1(_00945_),
    .C1(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__and2b_1 _08330_ (.A_N(_00939_),
    .B(_00941_),
    .X(_00948_));
 sky130_fd_sc_hd__o211a_1 _08331_ (.A1(_00946_),
    .A2(_00945_),
    .B1(_00944_),
    .C1(_00908_),
    .X(_00949_));
 sky130_fd_sc_hd__nor3_1 _08332_ (.A(_00947_),
    .B(_00948_),
    .C(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__or2_2 _08333_ (.A(_00947_),
    .B(_00950_),
    .X(_00951_));
 sky130_fd_sc_hd__a211oi_1 _08334_ (.A1(_00659_),
    .A2(_00660_),
    .B1(_00588_),
    .C1(_00621_),
    .Y(_00952_));
 sky130_fd_sc_hd__nor2_2 _08335_ (.A(_00661_),
    .B(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _08336_ (.A(_00951_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__a21oi_1 _08337_ (.A1(_00817_),
    .A2(_00818_),
    .B1(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__and3_1 _08338_ (.A(_00817_),
    .B(_00954_),
    .C(_00818_),
    .X(_00956_));
 sky130_fd_sc_hd__or3_1 _08339_ (.A(_00829_),
    .B(_00827_),
    .C(_00828_),
    .X(_00957_));
 sky130_fd_sc_hd__nand2_1 _08340_ (.A(_06460_),
    .B(_05241_),
    .Y(_00958_));
 sky130_fd_sc_hd__a22oi_2 _08341_ (.A1(_06463_),
    .A2(_05305_),
    .B1(_05370_),
    .B2(_06492_),
    .Y(_00959_));
 sky130_fd_sc_hd__and4_1 _08342_ (.A(_06469_),
    .B(_02194_),
    .C(net18),
    .D(net19),
    .X(_00960_));
 sky130_fd_sc_hd__o21bai_1 _08343_ (.A1(_00958_),
    .A2(_00959_),
    .B1_N(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__o21ai_1 _08344_ (.A1(_00829_),
    .A2(_00828_),
    .B1(_00827_),
    .Y(_00962_));
 sky130_fd_sc_hd__nand3_1 _08345_ (.A(_00957_),
    .B(_00961_),
    .C(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__a21o_1 _08346_ (.A1(_00957_),
    .A2(_00962_),
    .B1(_00961_),
    .X(_00964_));
 sky130_fd_sc_hd__nand2_1 _08347_ (.A(_06475_),
    .B(_00534_),
    .Y(_00965_));
 sky130_fd_sc_hd__a22oi_1 _08348_ (.A1(_06500_),
    .A2(_06517_),
    .B1(_06518_),
    .B2(_06501_),
    .Y(_00966_));
 sky130_fd_sc_hd__and4_1 _08349_ (.A(_06503_),
    .B(_06504_),
    .C(_05176_),
    .D(_05241_),
    .X(_00967_));
 sky130_fd_sc_hd__nor2_1 _08350_ (.A(_00966_),
    .B(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__xnor2_1 _08351_ (.A(_00965_),
    .B(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand3_1 _08352_ (.A(_00963_),
    .B(_00964_),
    .C(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__or3_1 _08353_ (.A(_00960_),
    .B(_00958_),
    .C(_00959_),
    .X(_00971_));
 sky130_fd_sc_hd__o21ai_1 _08354_ (.A1(_00960_),
    .A2(_00959_),
    .B1(_00958_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _08355_ (.A(_06488_),
    .B(_06517_),
    .Y(_00973_));
 sky130_fd_sc_hd__a22oi_2 _08356_ (.A1(_06491_),
    .A2(_05241_),
    .B1(_05305_),
    .B2(_06492_),
    .Y(_00974_));
 sky130_fd_sc_hd__and4_1 _08357_ (.A(_06494_),
    .B(_06495_),
    .C(_05241_),
    .D(_05305_),
    .X(_00975_));
 sky130_fd_sc_hd__o21bai_1 _08358_ (.A1(_00973_),
    .A2(_00974_),
    .B1_N(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__a21o_1 _08359_ (.A1(_00971_),
    .A2(_00972_),
    .B1(_00976_),
    .X(_00977_));
 sky130_fd_sc_hd__nand2_1 _08360_ (.A(net108),
    .B(_05025_),
    .Y(_00978_));
 sky130_fd_sc_hd__a22oi_1 _08361_ (.A1(_06504_),
    .A2(_05101_),
    .B1(_06517_),
    .B2(_06503_),
    .Y(_00979_));
 sky130_fd_sc_hd__and4_1 _08362_ (.A(net110),
    .B(net109),
    .C(net14),
    .D(_05176_),
    .X(_00980_));
 sky130_fd_sc_hd__nor2_1 _08363_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__xnor2_1 _08364_ (.A(_00978_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand3_1 _08365_ (.A(_00971_),
    .B(_00976_),
    .C(_00972_),
    .Y(_00983_));
 sky130_fd_sc_hd__a21bo_1 _08366_ (.A1(_00977_),
    .A2(_00982_),
    .B1_N(_00983_),
    .X(_00984_));
 sky130_fd_sc_hd__a21o_1 _08367_ (.A1(_00963_),
    .A2(_00964_),
    .B1(_00969_),
    .X(_00985_));
 sky130_fd_sc_hd__nand3_2 _08368_ (.A(_00970_),
    .B(_00984_),
    .C(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__a21o_1 _08369_ (.A1(_00970_),
    .A2(_00985_),
    .B1(_00984_),
    .X(_00987_));
 sky130_fd_sc_hd__and4_1 _08370_ (.A(_06519_),
    .B(net66),
    .C(net11),
    .D(net133),
    .X(_00988_));
 sky130_fd_sc_hd__nand2_1 _08371_ (.A(net106),
    .B(_06602_),
    .Y(_00989_));
 sky130_fd_sc_hd__a22oi_1 _08372_ (.A1(_02474_),
    .A2(_06604_),
    .B1(_06580_),
    .B2(_06564_),
    .Y(_00990_));
 sky130_fd_sc_hd__or3_1 _08373_ (.A(_00988_),
    .B(_00989_),
    .C(_00990_),
    .X(_00991_));
 sky130_fd_sc_hd__or2b_1 _08374_ (.A(_00988_),
    .B_N(_00991_),
    .X(_00992_));
 sky130_fd_sc_hd__and4_1 _08375_ (.A(net107),
    .B(net66),
    .C(net133),
    .D(net13),
    .X(_00993_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(net106),
    .B(_06604_),
    .Y(_00994_));
 sky130_fd_sc_hd__a22oi_2 _08377_ (.A1(_06515_),
    .A2(net133),
    .B1(_06581_),
    .B2(_06519_),
    .Y(_00995_));
 sky130_fd_sc_hd__or3_1 _08378_ (.A(_00993_),
    .B(_00994_),
    .C(_00995_),
    .X(_00996_));
 sky130_fd_sc_hd__o21bai_1 _08379_ (.A1(_00978_),
    .A2(_00979_),
    .B1_N(_00980_),
    .Y(_00997_));
 sky130_fd_sc_hd__o21ai_1 _08380_ (.A1(_00993_),
    .A2(_00995_),
    .B1(_00994_),
    .Y(_00998_));
 sky130_fd_sc_hd__and3_1 _08381_ (.A(_00996_),
    .B(_00997_),
    .C(_00998_),
    .X(_00999_));
 sky130_fd_sc_hd__a21o_1 _08382_ (.A1(_00996_),
    .A2(_00998_),
    .B1(_00997_),
    .X(_01000_));
 sky130_fd_sc_hd__and2b_1 _08383_ (.A_N(_00999_),
    .B(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__xor2_1 _08384_ (.A(_00992_),
    .B(_01001_),
    .X(_01002_));
 sky130_fd_sc_hd__nand3_1 _08385_ (.A(_00986_),
    .B(_00987_),
    .C(_01002_),
    .Y(_01003_));
 sky130_fd_sc_hd__nand3_1 _08386_ (.A(_00832_),
    .B(_00824_),
    .C(_00831_),
    .Y(_01004_));
 sky130_fd_sc_hd__a21bo_1 _08387_ (.A1(_00964_),
    .A2(_00969_),
    .B1_N(_00963_),
    .X(_01005_));
 sky130_fd_sc_hd__a21o_1 _08388_ (.A1(_00832_),
    .A2(_00831_),
    .B1(_00824_),
    .X(_01006_));
 sky130_fd_sc_hd__nand3_2 _08389_ (.A(_01004_),
    .B(_01005_),
    .C(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__a21o_1 _08390_ (.A1(_01004_),
    .A2(_01006_),
    .B1(_01005_),
    .X(_01008_));
 sky130_fd_sc_hd__and2b_1 _08391_ (.A_N(_00993_),
    .B(_00996_),
    .X(_01009_));
 sky130_fd_sc_hd__o21ba_1 _08392_ (.A1(_00965_),
    .A2(_00966_),
    .B1_N(_00967_),
    .X(_01010_));
 sky130_fd_sc_hd__nor2_1 _08393_ (.A(_00842_),
    .B(_00841_),
    .Y(_01011_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(_00840_),
    .B(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__xnor2_1 _08395_ (.A(_01010_),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__xnor2_1 _08396_ (.A(_01009_),
    .B(_01013_),
    .Y(_01014_));
 sky130_fd_sc_hd__a21oi_2 _08397_ (.A1(_01007_),
    .A2(_01008_),
    .B1(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _08398_ (.A(_01007_),
    .B(_01008_),
    .C(_01014_),
    .X(_01016_));
 sky130_fd_sc_hd__a211oi_4 _08399_ (.A1(_00986_),
    .A2(_01003_),
    .B1(_01015_),
    .C1(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__o211a_1 _08400_ (.A1(_01016_),
    .A2(_01015_),
    .B1(_01003_),
    .C1(_00986_),
    .X(_01018_));
 sky130_fd_sc_hd__and4_1 _08401_ (.A(_02593_),
    .B(_02658_),
    .C(_04778_),
    .D(_06603_),
    .X(_01019_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(_06593_),
    .B(_04714_),
    .Y(_01020_));
 sky130_fd_sc_hd__a22oi_2 _08403_ (.A1(_06682_),
    .A2(_06612_),
    .B1(_04843_),
    .B2(_00000_),
    .Y(_01021_));
 sky130_fd_sc_hd__or3_1 _08404_ (.A(_01019_),
    .B(_01020_),
    .C(_01021_),
    .X(_01022_));
 sky130_fd_sc_hd__o21ai_1 _08405_ (.A1(_01019_),
    .A2(_01021_),
    .B1(_01020_),
    .Y(_01023_));
 sky130_fd_sc_hd__a22o_1 _08406_ (.A1(_02647_),
    .A2(_00032_),
    .B1(_06611_),
    .B2(_02582_),
    .X(_01024_));
 sky130_fd_sc_hd__and4_1 _08407_ (.A(_02582_),
    .B(_02647_),
    .C(_00032_),
    .D(_04767_),
    .X(_01025_));
 sky130_fd_sc_hd__a31o_1 _08408_ (.A1(_02723_),
    .A2(_04660_),
    .A3(_01024_),
    .B1(_01025_),
    .X(_01026_));
 sky130_fd_sc_hd__nand3_1 _08409_ (.A(_01022_),
    .B(_01023_),
    .C(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21o_1 _08410_ (.A1(_01022_),
    .A2(_01023_),
    .B1(_01026_),
    .X(_01028_));
 sky130_fd_sc_hd__nand2_1 _08411_ (.A(_02851_),
    .B(_04531_),
    .Y(_01029_));
 sky130_fd_sc_hd__and4_1 _08412_ (.A(_06631_),
    .B(_06630_),
    .C(_04585_),
    .D(_00048_),
    .X(_01030_));
 sky130_fd_sc_hd__a22o_1 _08413_ (.A1(_06630_),
    .A2(_04585_),
    .B1(_04649_),
    .B2(_06631_),
    .X(_01031_));
 sky130_fd_sc_hd__and2b_1 _08414_ (.A_N(_01030_),
    .B(_01031_),
    .X(_01032_));
 sky130_fd_sc_hd__xnor2_2 _08415_ (.A(_01029_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand3_2 _08416_ (.A(_01027_),
    .B(_01028_),
    .C(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand2_1 _08417_ (.A(_01027_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__o21ai_1 _08418_ (.A1(_00852_),
    .A2(_00854_),
    .B1(_00853_),
    .Y(_01036_));
 sky130_fd_sc_hd__o21bai_1 _08419_ (.A1(_01020_),
    .A2(_01021_),
    .B1_N(_01019_),
    .Y(_01037_));
 sky130_fd_sc_hd__nand3_1 _08420_ (.A(_00855_),
    .B(_01036_),
    .C(_01037_),
    .Y(_01038_));
 sky130_fd_sc_hd__a21o_1 _08421_ (.A1(_00855_),
    .A2(_01036_),
    .B1(_01037_),
    .X(_01039_));
 sky130_fd_sc_hd__and3_1 _08422_ (.A(_00879_),
    .B(_00875_),
    .C(_00876_),
    .X(_01040_));
 sky130_fd_sc_hd__a21oi_1 _08423_ (.A1(_00879_),
    .A2(_00876_),
    .B1(_00875_),
    .Y(_01041_));
 sky130_fd_sc_hd__nor2_1 _08424_ (.A(_01040_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand3_1 _08425_ (.A(_01038_),
    .B(_01039_),
    .C(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__a21o_1 _08426_ (.A1(_00992_),
    .A2(_01000_),
    .B1(_00999_),
    .X(_01044_));
 sky130_fd_sc_hd__a21o_1 _08427_ (.A1(_01038_),
    .A2(_01039_),
    .B1(_01042_),
    .X(_01045_));
 sky130_fd_sc_hd__nand3_1 _08428_ (.A(_01043_),
    .B(_01044_),
    .C(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__a21o_1 _08429_ (.A1(_01043_),
    .A2(_01045_),
    .B1(_01044_),
    .X(_01047_));
 sky130_fd_sc_hd__nand3_1 _08430_ (.A(_01035_),
    .B(_01046_),
    .C(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__a21o_1 _08431_ (.A1(_01046_),
    .A2(_01047_),
    .B1(_01035_),
    .X(_01049_));
 sky130_fd_sc_hd__and4bb_1 _08432_ (.A_N(_01017_),
    .B_N(_01018_),
    .C(_01048_),
    .D(_01049_),
    .X(_01050_));
 sky130_fd_sc_hd__nand3_1 _08433_ (.A(_01007_),
    .B(_01008_),
    .C(_01014_),
    .Y(_01051_));
 sky130_fd_sc_hd__a21oi_1 _08434_ (.A1(_00835_),
    .A2(_00845_),
    .B1(_00844_),
    .Y(_01052_));
 sky130_fd_sc_hd__and3_1 _08435_ (.A(_00835_),
    .B(_00844_),
    .C(_00845_),
    .X(_01053_));
 sky130_fd_sc_hd__a211oi_1 _08436_ (.A1(_01007_),
    .A2(_01051_),
    .B1(_01052_),
    .C1(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__o211a_1 _08437_ (.A1(_01053_),
    .A2(_01052_),
    .B1(_01051_),
    .C1(_01007_),
    .X(_01055_));
 sky130_fd_sc_hd__nand2_1 _08438_ (.A(_01038_),
    .B(_01043_),
    .Y(_01056_));
 sky130_fd_sc_hd__or2b_1 _08439_ (.A(_01010_),
    .B_N(_01012_),
    .X(_01057_));
 sky130_fd_sc_hd__or2b_1 _08440_ (.A(_01009_),
    .B_N(_01013_),
    .X(_01058_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(_00858_),
    .B(_00861_),
    .Y(_01059_));
 sky130_fd_sc_hd__a21o_1 _08442_ (.A1(_01057_),
    .A2(_01058_),
    .B1(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__nand3_1 _08443_ (.A(_01057_),
    .B(_01058_),
    .C(_01059_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand3_2 _08444_ (.A(_01056_),
    .B(_01060_),
    .C(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__a21o_1 _08445_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_01056_),
    .X(_01063_));
 sky130_fd_sc_hd__a2bb2o_1 _08446_ (.A1_N(_01054_),
    .A2_N(_01055_),
    .B1(_01062_),
    .B2(_01063_),
    .X(_01064_));
 sky130_fd_sc_hd__or4bb_4 _08447_ (.A(_01054_),
    .B(_01055_),
    .C_N(_01062_),
    .D_N(_01063_),
    .X(_01065_));
 sky130_fd_sc_hd__o211ai_4 _08448_ (.A1(_01017_),
    .A2(_01050_),
    .B1(_01064_),
    .C1(_01065_),
    .Y(_01066_));
 sky130_fd_sc_hd__a211o_1 _08449_ (.A1(_01065_),
    .A2(_01064_),
    .B1(_01050_),
    .C1(_01017_),
    .X(_01067_));
 sky130_fd_sc_hd__a31o_1 _08450_ (.A1(_02840_),
    .A2(_04531_),
    .A3(_01031_),
    .B1(_01030_),
    .X(_01068_));
 sky130_fd_sc_hd__o21ai_1 _08451_ (.A1(_00883_),
    .A2(_00885_),
    .B1(_00884_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand3_1 _08452_ (.A(_00886_),
    .B(_01068_),
    .C(_01069_),
    .Y(_01070_));
 sky130_fd_sc_hd__and4_1 _08453_ (.A(net120),
    .B(net44),
    .C(_00089_),
    .D(_00082_),
    .X(_01071_));
 sky130_fd_sc_hd__nand2_1 _08454_ (.A(net119),
    .B(_04294_),
    .Y(_01072_));
 sky130_fd_sc_hd__a22oi_2 _08455_ (.A1(_00029_),
    .A2(_00072_),
    .B1(_00083_),
    .B2(_00028_),
    .Y(_01073_));
 sky130_fd_sc_hd__or3_1 _08456_ (.A(_01071_),
    .B(_01072_),
    .C(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__or2b_1 _08457_ (.A(_01071_),
    .B_N(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__a21o_1 _08458_ (.A1(_00886_),
    .A2(_01069_),
    .B1(_01068_),
    .X(_01076_));
 sky130_fd_sc_hd__nand3_1 _08459_ (.A(_01070_),
    .B(_01075_),
    .C(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__a21o_1 _08460_ (.A1(_01070_),
    .A2(_01076_),
    .B1(_01075_),
    .X(_01078_));
 sky130_fd_sc_hd__and4_1 _08461_ (.A(_00028_),
    .B(_00029_),
    .C(_04294_),
    .D(_00072_),
    .X(_01079_));
 sky130_fd_sc_hd__a22oi_1 _08462_ (.A1(_00046_),
    .A2(_00074_),
    .B1(_00090_),
    .B2(_00049_),
    .Y(_01080_));
 sky130_fd_sc_hd__nor2_1 _08463_ (.A(_01079_),
    .B(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__a31o_1 _08464_ (.A1(_00221_),
    .A2(_04251_),
    .A3(_01081_),
    .B1(_01079_),
    .X(_01082_));
 sky130_fd_sc_hd__o21ai_1 _08465_ (.A1(_01071_),
    .A2(_01073_),
    .B1(_01072_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _08466_ (.A(net121),
    .B(_04445_),
    .Y(_01084_));
 sky130_fd_sc_hd__a22oi_1 _08467_ (.A1(_06601_),
    .A2(_00085_),
    .B1(_04585_),
    .B2(_06606_),
    .Y(_01085_));
 sky130_fd_sc_hd__and4_1 _08468_ (.A(_06598_),
    .B(_06599_),
    .C(_04509_),
    .D(_00035_),
    .X(_01086_));
 sky130_fd_sc_hd__o21bai_1 _08469_ (.A1(_01084_),
    .A2(_01085_),
    .B1_N(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__a21o_1 _08470_ (.A1(_01074_),
    .A2(_01083_),
    .B1(_01087_),
    .X(_01088_));
 sky130_fd_sc_hd__nand3_1 _08471_ (.A(_01074_),
    .B(_01087_),
    .C(_01083_),
    .Y(_01089_));
 sky130_fd_sc_hd__a21bo_1 _08472_ (.A1(_01082_),
    .A2(_01088_),
    .B1_N(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__and3_1 _08473_ (.A(_01077_),
    .B(_01078_),
    .C(_01090_),
    .X(_01091_));
 sky130_fd_sc_hd__inv_2 _08474_ (.A(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21oi_1 _08475_ (.A1(_01077_),
    .A2(_01078_),
    .B1(_01090_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(_03335_),
    .B(_03982_),
    .Y(_01094_));
 sky130_fd_sc_hd__and2b_1 _08477_ (.A_N(_00913_),
    .B(_00912_),
    .X(_01095_));
 sky130_fd_sc_hd__xnor2_2 _08478_ (.A(_01094_),
    .B(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_1 _08479_ (.A(_00923_),
    .B(_00922_),
    .Y(_01097_));
 sky130_fd_sc_hd__xnor2_1 _08480_ (.A(_00920_),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__and4_1 _08481_ (.A(_00095_),
    .B(_00096_),
    .C(_00271_),
    .D(_04229_),
    .X(_01099_));
 sky130_fd_sc_hd__a22oi_1 _08482_ (.A1(_03099_),
    .A2(_04176_),
    .B1(_04240_),
    .B2(_03056_),
    .Y(_01100_));
 sky130_fd_sc_hd__and4bb_1 _08483_ (.A_N(_01099_),
    .B_N(_01100_),
    .C(_03163_),
    .D(_00303_),
    .X(_01101_));
 sky130_fd_sc_hd__nor2_2 _08484_ (.A(_01099_),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__xnor2_1 _08485_ (.A(_01098_),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__xnor2_1 _08486_ (.A(_01096_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__or3_1 _08487_ (.A(_01091_),
    .B(_01093_),
    .C(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__a21o_1 _08488_ (.A1(_00882_),
    .A2(_00888_),
    .B1(_00887_),
    .X(_01106_));
 sky130_fd_sc_hd__a21bo_1 _08489_ (.A1(_01075_),
    .A2(_01076_),
    .B1_N(_01070_),
    .X(_01107_));
 sky130_fd_sc_hd__and3_1 _08490_ (.A(_00889_),
    .B(_01106_),
    .C(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__a21oi_1 _08491_ (.A1(_00889_),
    .A2(_01106_),
    .B1(_01107_),
    .Y(_01109_));
 sky130_fd_sc_hd__and2b_1 _08492_ (.A_N(_00926_),
    .B(_00925_),
    .X(_01110_));
 sky130_fd_sc_hd__xnor2_1 _08493_ (.A(_00918_),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__o21a_1 _08494_ (.A1(_01108_),
    .A2(_01109_),
    .B1(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__nor3_1 _08495_ (.A(_01108_),
    .B(_01109_),
    .C(_01111_),
    .Y(_01113_));
 sky130_fd_sc_hd__a211oi_2 _08496_ (.A1(_01046_),
    .A2(_01048_),
    .B1(_01112_),
    .C1(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__o211a_1 _08497_ (.A1(_01113_),
    .A2(_01112_),
    .B1(_01048_),
    .C1(_01046_),
    .X(_01115_));
 sky130_fd_sc_hd__a211oi_1 _08498_ (.A1(_01092_),
    .A2(_01105_),
    .B1(_01114_),
    .C1(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__inv_2 _08499_ (.A(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hd__o211ai_2 _08500_ (.A1(_01114_),
    .A2(_01115_),
    .B1(_01092_),
    .C1(_01105_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand4_1 _08501_ (.A(_01066_),
    .B(_01067_),
    .C(_01117_),
    .D(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__a211o_1 _08502_ (.A1(_01007_),
    .A2(_01051_),
    .B1(_01052_),
    .C1(_01053_),
    .X(_01120_));
 sky130_fd_sc_hd__o211a_1 _08503_ (.A1(_00848_),
    .A2(_00847_),
    .B1(_00846_),
    .C1(_00835_),
    .X(_01121_));
 sky130_fd_sc_hd__o2bb2a_1 _08504_ (.A1_N(_00868_),
    .A2_N(_00869_),
    .B1(_01121_),
    .B2(_00849_),
    .X(_01122_));
 sky130_fd_sc_hd__a211oi_1 _08505_ (.A1(_01120_),
    .A2(_01065_),
    .B1(_01122_),
    .C1(_00871_),
    .Y(_01123_));
 sky130_fd_sc_hd__o211a_1 _08506_ (.A1(_00871_),
    .A2(_01122_),
    .B1(_01065_),
    .C1(_01120_),
    .X(_01124_));
 sky130_fd_sc_hd__inv_2 _08507_ (.A(_01108_),
    .Y(_01125_));
 sky130_fd_sc_hd__or3_1 _08508_ (.A(_01108_),
    .B(_01109_),
    .C(_01111_),
    .X(_01126_));
 sky130_fd_sc_hd__o21a_1 _08509_ (.A1(_00892_),
    .A2(_00893_),
    .B1(_00896_),
    .X(_01127_));
 sky130_fd_sc_hd__nor3_2 _08510_ (.A(_00892_),
    .B(_00893_),
    .C(_00896_),
    .Y(_01128_));
 sky130_fd_sc_hd__a211oi_4 _08511_ (.A1(_01060_),
    .A2(_01062_),
    .B1(_01127_),
    .C1(_01128_),
    .Y(_01129_));
 sky130_fd_sc_hd__o211a_1 _08512_ (.A1(_01128_),
    .A2(_01127_),
    .B1(_01062_),
    .C1(_01060_),
    .X(_01130_));
 sky130_fd_sc_hd__a211oi_4 _08513_ (.A1(_01125_),
    .A2(_01126_),
    .B1(_01129_),
    .C1(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__o211a_1 _08514_ (.A1(_01129_),
    .A2(_01130_),
    .B1(_01125_),
    .C1(_01126_),
    .X(_01132_));
 sky130_fd_sc_hd__o22a_1 _08515_ (.A1(_01123_),
    .A2(_01124_),
    .B1(_01131_),
    .B2(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__nor4_2 _08516_ (.A(_01123_),
    .B(_01124_),
    .C(_01131_),
    .D(_01132_),
    .Y(_01134_));
 sky130_fd_sc_hd__a211oi_2 _08517_ (.A1(_01066_),
    .A2(_01119_),
    .B1(_01133_),
    .C1(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__o211a_1 _08518_ (.A1(_01134_),
    .A2(_01133_),
    .B1(_01119_),
    .C1(_01066_),
    .X(_01136_));
 sky130_fd_sc_hd__nor2_1 _08519_ (.A(_01114_),
    .B(_01116_),
    .Y(_01137_));
 sky130_fd_sc_hd__and2b_1 _08520_ (.A_N(_01102_),
    .B(_01098_),
    .X(_01138_));
 sky130_fd_sc_hd__and2_1 _08521_ (.A(_01096_),
    .B(_01103_),
    .X(_01139_));
 sky130_fd_sc_hd__and2b_1 _08522_ (.A_N(_00914_),
    .B(_00911_),
    .X(_01140_));
 sky130_fd_sc_hd__nor2_1 _08523_ (.A(_00915_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__o21ai_1 _08524_ (.A1(_01138_),
    .A2(_01139_),
    .B1(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__or3_1 _08525_ (.A(_01138_),
    .B(_01139_),
    .C(_01141_),
    .X(_01143_));
 sky130_fd_sc_hd__and4_1 _08526_ (.A(_03217_),
    .B(_03271_),
    .C(net132),
    .D(_06430_),
    .X(_01144_));
 sky130_fd_sc_hd__inv_2 _08527_ (.A(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__buf_4 _08528_ (.A(_03271_),
    .X(_01146_));
 sky130_fd_sc_hd__clkbuf_8 _08529_ (.A(_03217_),
    .X(_01147_));
 sky130_fd_sc_hd__a22o_1 _08530_ (.A1(_01146_),
    .A2(_06437_),
    .B1(_06443_),
    .B2(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__and4_1 _08531_ (.A(_03335_),
    .B(_03884_),
    .C(_01145_),
    .D(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__o211a_1 _08532_ (.A1(_01144_),
    .A2(_01149_),
    .B1(_03400_),
    .C1(_03906_),
    .X(_01150_));
 sky130_fd_sc_hd__nand2_1 _08533_ (.A(_01143_),
    .B(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__xnor2_1 _08534_ (.A(_00915_),
    .B(_00930_),
    .Y(_01152_));
 sky130_fd_sc_hd__a21o_1 _08535_ (.A1(_01142_),
    .A2(_01151_),
    .B1(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__nand3_1 _08536_ (.A(_01152_),
    .B(_01142_),
    .C(_01151_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _08537_ (.A(_01153_),
    .B(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__xnor2_1 _08538_ (.A(_01137_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__and2_1 _08539_ (.A(_01143_),
    .B(_01142_),
    .X(_01157_));
 sky130_fd_sc_hd__and4_1 _08540_ (.A(_00237_),
    .B(_00462_),
    .C(_06431_),
    .D(_00287_),
    .X(_01158_));
 sky130_fd_sc_hd__a22oi_1 _08541_ (.A1(_00132_),
    .A2(_06433_),
    .B1(_04176_),
    .B2(_00133_),
    .Y(_01159_));
 sky130_fd_sc_hd__and4bb_1 _08542_ (.A_N(_01158_),
    .B_N(_01159_),
    .C(_03163_),
    .D(_06443_),
    .X(_01160_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_01158_),
    .B(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__o2bb2a_1 _08544_ (.A1_N(_00262_),
    .A2_N(_00303_),
    .B1(_01099_),
    .B2(_01100_),
    .X(_01162_));
 sky130_fd_sc_hd__nor2_1 _08545_ (.A(_01101_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__and2b_1 _08546_ (.A_N(_01161_),
    .B(_01163_),
    .X(_01164_));
 sky130_fd_sc_hd__a22oi_1 _08547_ (.A1(_03335_),
    .A2(_03884_),
    .B1(_01145_),
    .B2(_01148_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _08548_ (.A(_01149_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_01163_),
    .B(_01161_),
    .Y(_01167_));
 sky130_fd_sc_hd__and2_1 _08550_ (.A(_01166_),
    .B(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__a211oi_1 _08551_ (.A1(_03400_),
    .A2(_03906_),
    .B1(_01144_),
    .C1(_01149_),
    .Y(_01169_));
 sky130_fd_sc_hd__or2_1 _08552_ (.A(_01150_),
    .B(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__o21ba_1 _08553_ (.A1(_01164_),
    .A2(_01168_),
    .B1_N(_01170_),
    .X(_01171_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_01157_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__xnor2_1 _08555_ (.A(_01156_),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor3_1 _08556_ (.A(_01135_),
    .B(_01136_),
    .C(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__and4_1 _08557_ (.A(_00874_),
    .B(_00902_),
    .C(_00903_),
    .D(_00904_),
    .X(_01175_));
 sky130_fd_sc_hd__a211o_1 _08558_ (.A1(_01120_),
    .A2(_01065_),
    .B1(_01122_),
    .C1(_00871_),
    .X(_01176_));
 sky130_fd_sc_hd__o31a_1 _08559_ (.A1(_01124_),
    .A2(_01131_),
    .A3(_01132_),
    .B1(_01176_),
    .X(_01177_));
 sky130_fd_sc_hd__a22oi_2 _08560_ (.A1(_00902_),
    .A2(_00903_),
    .B1(_00904_),
    .B2(_00874_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor3_1 _08561_ (.A(_01175_),
    .B(_01177_),
    .C(_01178_),
    .Y(_01179_));
 sky130_fd_sc_hd__o21a_1 _08562_ (.A1(_01175_),
    .A2(_01178_),
    .B1(_01177_),
    .X(_01180_));
 sky130_fd_sc_hd__xor2_1 _08563_ (.A(_00934_),
    .B(_00935_),
    .X(_01181_));
 sky130_fd_sc_hd__o21a_1 _08564_ (.A1(_01129_),
    .A2(_01131_),
    .B1(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__nor3_1 _08565_ (.A(_01129_),
    .B(_01131_),
    .C(_01181_),
    .Y(_01183_));
 sky130_fd_sc_hd__nor3_2 _08566_ (.A(_01153_),
    .B(_01182_),
    .C(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__o21a_1 _08567_ (.A1(_01182_),
    .A2(_01183_),
    .B1(_01153_),
    .X(_01185_));
 sky130_fd_sc_hd__o22ai_2 _08568_ (.A1(_01179_),
    .A2(_01180_),
    .B1(_01184_),
    .B2(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__or4_2 _08569_ (.A(_01179_),
    .B(_01180_),
    .C(_01184_),
    .D(_01185_),
    .X(_01187_));
 sky130_fd_sc_hd__o211a_2 _08570_ (.A1(_01135_),
    .A2(_01174_),
    .B1(_01186_),
    .C1(_01187_),
    .X(_01188_));
 sky130_fd_sc_hd__or2_1 _08571_ (.A(_01156_),
    .B(_01172_),
    .X(_01189_));
 sky130_fd_sc_hd__o21a_1 _08572_ (.A1(_01137_),
    .A2(_01155_),
    .B1(_01189_),
    .X(_01190_));
 sky130_fd_sc_hd__a211oi_1 _08573_ (.A1(_01187_),
    .A2(_01186_),
    .B1(_01174_),
    .C1(_01135_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor3_1 _08574_ (.A(_01188_),
    .B(_01190_),
    .C(_01191_),
    .Y(_01192_));
 sky130_fd_sc_hd__or3_1 _08575_ (.A(_01175_),
    .B(_01177_),
    .C(_01178_),
    .X(_01193_));
 sky130_fd_sc_hd__a22oi_2 _08576_ (.A1(_00941_),
    .A2(_00942_),
    .B1(_00943_),
    .B2(_00908_),
    .Y(_01194_));
 sky130_fd_sc_hd__and4_1 _08577_ (.A(_00908_),
    .B(_00941_),
    .C(_00942_),
    .D(_00943_),
    .X(_01195_));
 sky130_fd_sc_hd__a211o_2 _08578_ (.A1(_01193_),
    .A2(_01187_),
    .B1(_01194_),
    .C1(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__o211ai_2 _08579_ (.A1(_01195_),
    .A2(_01194_),
    .B1(_01187_),
    .C1(_01193_),
    .Y(_01197_));
 sky130_fd_sc_hd__a211o_1 _08580_ (.A1(_01196_),
    .A2(_01197_),
    .B1(_01182_),
    .C1(_01184_),
    .X(_01198_));
 sky130_fd_sc_hd__o211ai_4 _08581_ (.A1(_01182_),
    .A2(_01184_),
    .B1(_01196_),
    .C1(_01197_),
    .Y(_01199_));
 sky130_fd_sc_hd__o211ai_4 _08582_ (.A1(_01188_),
    .A2(_01192_),
    .B1(_01198_),
    .C1(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__a211o_1 _08583_ (.A1(_01199_),
    .A2(_01198_),
    .B1(_01192_),
    .C1(_01188_),
    .X(_01201_));
 sky130_fd_sc_hd__or3_1 _08584_ (.A(_01188_),
    .B(_01190_),
    .C(_01191_),
    .X(_01202_));
 sky130_fd_sc_hd__and4_1 _08585_ (.A(_03239_),
    .B(_03293_),
    .C(_03884_),
    .D(_03982_),
    .X(_01203_));
 sky130_fd_sc_hd__and4_1 _08586_ (.A(_00095_),
    .B(_00096_),
    .C(_06430_),
    .D(_06431_),
    .X(_01204_));
 sky130_fd_sc_hd__inv_2 _08587_ (.A(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__buf_4 _08588_ (.A(_00462_),
    .X(_01206_));
 sky130_fd_sc_hd__a22o_1 _08589_ (.A1(_01206_),
    .A2(_06446_),
    .B1(_00303_),
    .B2(_00921_),
    .X(_01207_));
 sky130_fd_sc_hd__and4_1 _08590_ (.A(_03174_),
    .B(_03971_),
    .C(_01205_),
    .D(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__o2bb2a_1 _08591_ (.A1_N(_03174_),
    .A2_N(_04057_),
    .B1(_01158_),
    .B2(_01159_),
    .X(_01209_));
 sky130_fd_sc_hd__nor2_2 _08592_ (.A(_01160_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__o21a_1 _08593_ (.A1(_01204_),
    .A2(_01208_),
    .B1(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__or3b_1 _08594_ (.A(_01164_),
    .B(_01168_),
    .C_N(_01170_),
    .X(_01212_));
 sky130_fd_sc_hd__and2b_1 _08595_ (.A_N(_01171_),
    .B(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__and3_1 _08596_ (.A(_01203_),
    .B(_01211_),
    .C(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__and4_1 _08597_ (.A(_02420_),
    .B(_06513_),
    .C(_06602_),
    .D(_06604_),
    .X(_01215_));
 sky130_fd_sc_hd__a22oi_1 _08598_ (.A1(_02485_),
    .A2(_04832_),
    .B1(_04896_),
    .B2(_06565_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _08599_ (.A(_01215_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__a31o_1 _08600_ (.A1(_02539_),
    .A2(_06613_),
    .A3(_01217_),
    .B1(_01215_),
    .X(_01218_));
 sky130_fd_sc_hd__o21ai_1 _08601_ (.A1(_00988_),
    .A2(_00990_),
    .B1(_00989_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(net108),
    .B(_04961_),
    .Y(_01220_));
 sky130_fd_sc_hd__a22oi_1 _08603_ (.A1(_06500_),
    .A2(_05025_),
    .B1(_06623_),
    .B2(_06501_),
    .Y(_01221_));
 sky130_fd_sc_hd__and4_1 _08604_ (.A(_06479_),
    .B(_06480_),
    .C(_06581_),
    .D(_05101_),
    .X(_01222_));
 sky130_fd_sc_hd__o21bai_1 _08605_ (.A1(_01220_),
    .A2(_01221_),
    .B1_N(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__a21o_1 _08606_ (.A1(_00991_),
    .A2(_01219_),
    .B1(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__and3_1 _08607_ (.A(_00991_),
    .B(_01223_),
    .C(_01219_),
    .X(_01225_));
 sky130_fd_sc_hd__a21o_1 _08608_ (.A1(_01218_),
    .A2(_01224_),
    .B1(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__a21o_1 _08609_ (.A1(_01027_),
    .A2(_01028_),
    .B1(_01033_),
    .X(_01227_));
 sky130_fd_sc_hd__nand3_4 _08610_ (.A(_01034_),
    .B(_01226_),
    .C(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__and4_1 _08611_ (.A(_06578_),
    .B(_06579_),
    .C(_00030_),
    .D(_04703_),
    .X(_01229_));
 sky130_fd_sc_hd__a22oi_1 _08612_ (.A1(_06583_),
    .A2(_04638_),
    .B1(_00033_),
    .B2(_06585_),
    .Y(_01230_));
 sky130_fd_sc_hd__and4bb_1 _08613_ (.A_N(_01229_),
    .B_N(_01230_),
    .C(_02712_),
    .D(_04585_),
    .X(_01231_));
 sky130_fd_sc_hd__nor2_1 _08614_ (.A(_01229_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_2 _08615_ (.A(_06593_),
    .B(_04649_),
    .Y(_01233_));
 sky130_fd_sc_hd__and2b_1 _08616_ (.A_N(_01025_),
    .B(_01024_),
    .X(_01234_));
 sky130_fd_sc_hd__xnor2_2 _08617_ (.A(_01233_),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__and2b_1 _08618_ (.A_N(_01232_),
    .B(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_1 _08619_ (.A(_01235_),
    .B(_01232_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _08620_ (.A(_01086_),
    .B(_01085_),
    .Y(_01238_));
 sky130_fd_sc_hd__xnor2_1 _08621_ (.A(_01084_),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__and2_1 _08622_ (.A(_01237_),
    .B(_01239_),
    .X(_01240_));
 sky130_fd_sc_hd__a21o_1 _08623_ (.A1(_01034_),
    .A2(_01227_),
    .B1(_01226_),
    .X(_01241_));
 sky130_fd_sc_hd__o211ai_4 _08624_ (.A1(_01236_),
    .A2(_01240_),
    .B1(_01228_),
    .C1(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__o21a_1 _08625_ (.A1(_01091_),
    .A2(_01093_),
    .B1(_01104_),
    .X(_01243_));
 sky130_fd_sc_hd__nor3_2 _08626_ (.A(_01091_),
    .B(_01093_),
    .C(_01104_),
    .Y(_01244_));
 sky130_fd_sc_hd__a211oi_4 _08627_ (.A1(_01228_),
    .A2(_01242_),
    .B1(_01243_),
    .C1(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__and4_1 _08628_ (.A(_02754_),
    .B(_02797_),
    .C(_00083_),
    .D(_00098_),
    .X(_01246_));
 sky130_fd_sc_hd__a22oi_1 _08629_ (.A1(_06601_),
    .A2(_04445_),
    .B1(_00085_),
    .B2(_06606_),
    .Y(_01247_));
 sky130_fd_sc_hd__and4bb_1 _08630_ (.A_N(_01246_),
    .B_N(_01247_),
    .C(_06608_),
    .D(_04369_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _08631_ (.A(_01246_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_00444_),
    .B(_00301_),
    .Y(_01250_));
 sky130_fd_sc_hd__xnor2_2 _08633_ (.A(_01250_),
    .B(_01081_),
    .Y(_01251_));
 sky130_fd_sc_hd__or2b_1 _08634_ (.A(_01249_),
    .B_N(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__and4_1 _08635_ (.A(_02894_),
    .B(_02948_),
    .C(_00267_),
    .D(_00074_),
    .X(_01253_));
 sky130_fd_sc_hd__a22oi_1 _08636_ (.A1(_00062_),
    .A2(_04240_),
    .B1(_04305_),
    .B2(_00063_),
    .Y(_01254_));
 sky130_fd_sc_hd__and4bb_1 _08637_ (.A_N(_01253_),
    .B_N(_01254_),
    .C(_03002_),
    .D(_00272_),
    .X(_01255_));
 sky130_fd_sc_hd__or2_1 _08638_ (.A(_01253_),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__xnor2_1 _08639_ (.A(_01249_),
    .B(_01251_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _08640_ (.A(_01256_),
    .B(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__and3_1 _08641_ (.A(_01089_),
    .B(_01082_),
    .C(_01088_),
    .X(_01259_));
 sky130_fd_sc_hd__a21oi_1 _08642_ (.A1(_01089_),
    .A2(_01088_),
    .B1(_01082_),
    .Y(_01260_));
 sky130_fd_sc_hd__or2_1 _08643_ (.A(_01259_),
    .B(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__a21oi_2 _08644_ (.A1(_01252_),
    .A2(_01258_),
    .B1(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__inv_2 _08645_ (.A(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__and3_1 _08646_ (.A(_01261_),
    .B(_01252_),
    .C(_01258_),
    .X(_01264_));
 sky130_fd_sc_hd__nor2_1 _08647_ (.A(_01166_),
    .B(_01167_),
    .Y(_01265_));
 sky130_fd_sc_hd__or2_2 _08648_ (.A(_01168_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__or3_2 _08649_ (.A(_01262_),
    .B(_01264_),
    .C(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__o211a_1 _08650_ (.A1(_01244_),
    .A2(_01243_),
    .B1(_01242_),
    .C1(_01228_),
    .X(_01268_));
 sky130_fd_sc_hd__a211oi_2 _08651_ (.A1(_01263_),
    .A2(_01267_),
    .B1(_01245_),
    .C1(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _08652_ (.A(_01150_),
    .B(_01171_),
    .Y(_01270_));
 sky130_fd_sc_hd__xnor2_1 _08653_ (.A(_01157_),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__o21a_1 _08654_ (.A1(_01245_),
    .A2(_01269_),
    .B1(_01271_),
    .X(_01272_));
 sky130_fd_sc_hd__nor3_1 _08655_ (.A(_01245_),
    .B(_01269_),
    .C(_01271_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _08656_ (.A(_01272_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__a21o_1 _08657_ (.A1(_01214_),
    .A2(_01274_),
    .B1(_01272_),
    .X(_01275_));
 sky130_fd_sc_hd__or3_1 _08658_ (.A(_01135_),
    .B(_01136_),
    .C(_01173_),
    .X(_01276_));
 sky130_fd_sc_hd__o21ai_1 _08659_ (.A1(_01135_),
    .A2(_01136_),
    .B1(_01173_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand3_1 _08660_ (.A(_00983_),
    .B(_00977_),
    .C(_00982_),
    .Y(_01278_));
 sky130_fd_sc_hd__or3_1 _08661_ (.A(_00975_),
    .B(_00973_),
    .C(_00974_),
    .X(_01279_));
 sky130_fd_sc_hd__o21ai_1 _08662_ (.A1(_00975_),
    .A2(_00974_),
    .B1(_00973_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _08663_ (.A(_06460_),
    .B(_05101_),
    .Y(_01281_));
 sky130_fd_sc_hd__a22oi_2 _08664_ (.A1(_06495_),
    .A2(_05176_),
    .B1(_05241_),
    .B2(_02107_),
    .Y(_01282_));
 sky130_fd_sc_hd__and4_1 _08665_ (.A(_02096_),
    .B(_02194_),
    .C(_05176_),
    .D(net17),
    .X(_01283_));
 sky130_fd_sc_hd__o21bai_1 _08666_ (.A1(_01281_),
    .A2(_01282_),
    .B1_N(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__a21o_1 _08667_ (.A1(_01279_),
    .A2(_01280_),
    .B1(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__nor2_1 _08668_ (.A(_01221_),
    .B(_01222_),
    .Y(_01286_));
 sky130_fd_sc_hd__xnor2_1 _08669_ (.A(_01220_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand3_1 _08670_ (.A(_01279_),
    .B(_01284_),
    .C(_01280_),
    .Y(_01288_));
 sky130_fd_sc_hd__a21bo_1 _08671_ (.A1(_01285_),
    .A2(_01287_),
    .B1_N(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__a21o_1 _08672_ (.A1(_00983_),
    .A2(_00977_),
    .B1(_00982_),
    .X(_01290_));
 sky130_fd_sc_hd__nand3_2 _08673_ (.A(_01278_),
    .B(_01289_),
    .C(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__a21o_1 _08674_ (.A1(_01278_),
    .A2(_01290_),
    .B1(_01289_),
    .X(_01292_));
 sky130_fd_sc_hd__and2b_1 _08675_ (.A_N(_01225_),
    .B(_01224_),
    .X(_01293_));
 sky130_fd_sc_hd__xor2_1 _08676_ (.A(_01218_),
    .B(_01293_),
    .X(_01294_));
 sky130_fd_sc_hd__nand3_1 _08677_ (.A(_01291_),
    .B(_01292_),
    .C(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__a21oi_2 _08678_ (.A1(_00986_),
    .A2(_00987_),
    .B1(_01002_),
    .Y(_01296_));
 sky130_fd_sc_hd__and3_1 _08679_ (.A(_00986_),
    .B(_00987_),
    .C(_01002_),
    .X(_01297_));
 sky130_fd_sc_hd__a211oi_4 _08680_ (.A1(_01291_),
    .A2(_01295_),
    .B1(_01296_),
    .C1(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__o211a_1 _08681_ (.A1(_01297_),
    .A2(_01296_),
    .B1(_01295_),
    .C1(_01291_),
    .X(_01299_));
 sky130_fd_sc_hd__a211o_1 _08682_ (.A1(_01228_),
    .A2(_01241_),
    .B1(_01236_),
    .C1(_01240_),
    .X(_01300_));
 sky130_fd_sc_hd__and4bb_1 _08683_ (.A_N(_01298_),
    .B_N(_01299_),
    .C(_01242_),
    .D(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__a2bb2o_1 _08684_ (.A1_N(_01017_),
    .A2_N(_01018_),
    .B1(_01048_),
    .B2(_01049_),
    .X(_01302_));
 sky130_fd_sc_hd__or4bb_2 _08685_ (.A(_01017_),
    .B(_01018_),
    .C_N(_01048_),
    .D_N(_01049_),
    .X(_01303_));
 sky130_fd_sc_hd__o211ai_4 _08686_ (.A1(_01298_),
    .A2(_01301_),
    .B1(_01302_),
    .C1(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__a211o_1 _08687_ (.A1(_01303_),
    .A2(_01302_),
    .B1(_01301_),
    .C1(_01298_),
    .X(_01305_));
 sky130_fd_sc_hd__inv_2 _08688_ (.A(_01269_),
    .Y(_01306_));
 sky130_fd_sc_hd__o211ai_4 _08689_ (.A1(_01245_),
    .A2(_01268_),
    .B1(_01263_),
    .C1(_01267_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand4_1 _08690_ (.A(_01304_),
    .B(_01305_),
    .C(_01306_),
    .D(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__a22oi_2 _08691_ (.A1(_01066_),
    .A2(_01067_),
    .B1(_01117_),
    .B2(_01118_),
    .Y(_01309_));
 sky130_fd_sc_hd__and4_1 _08692_ (.A(_01066_),
    .B(_01067_),
    .C(_01117_),
    .D(_01118_),
    .X(_01310_));
 sky130_fd_sc_hd__a211oi_2 _08693_ (.A1(_01304_),
    .A2(_01308_),
    .B1(_01309_),
    .C1(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__o211a_1 _08694_ (.A1(_01310_),
    .A2(_01309_),
    .B1(_01308_),
    .C1(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__xnor2_1 _08695_ (.A(_01214_),
    .B(_01274_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor3_1 _08696_ (.A(_01311_),
    .B(_01312_),
    .C(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__a211o_1 _08697_ (.A1(_01276_),
    .A2(_01277_),
    .B1(_01314_),
    .C1(_01311_),
    .X(_01315_));
 sky130_fd_sc_hd__o211ai_1 _08698_ (.A1(_01311_),
    .A2(_01314_),
    .B1(_01277_),
    .C1(_01276_),
    .Y(_01316_));
 sky130_fd_sc_hd__a21bo_1 _08699_ (.A1(_01275_),
    .A2(_01315_),
    .B1_N(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__o21ai_1 _08700_ (.A1(_01188_),
    .A2(_01191_),
    .B1(_01190_),
    .Y(_01318_));
 sky130_fd_sc_hd__and3_1 _08701_ (.A(_01202_),
    .B(_01317_),
    .C(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__nand3_1 _08702_ (.A(_01200_),
    .B(_01201_),
    .C(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__a21o_1 _08703_ (.A1(_01200_),
    .A2(_01201_),
    .B1(_01319_),
    .X(_01321_));
 sky130_fd_sc_hd__and2_1 _08704_ (.A(_01320_),
    .B(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__nand2_2 _08705_ (.A(_01196_),
    .B(_01199_),
    .Y(_01323_));
 sky130_fd_sc_hd__o21a_1 _08706_ (.A1(_00947_),
    .A2(_00949_),
    .B1(_00948_),
    .X(_01324_));
 sky130_fd_sc_hd__nor2_2 _08707_ (.A(_00950_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__xnor2_2 _08708_ (.A(_01323_),
    .B(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__xor2_4 _08709_ (.A(_01200_),
    .B(_01326_),
    .X(_01327_));
 sky130_fd_sc_hd__xnor2_2 _08710_ (.A(_00951_),
    .B(_00953_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _08711_ (.A(_01323_),
    .B(_01325_),
    .Y(_01329_));
 sky130_fd_sc_hd__xor2_2 _08712_ (.A(_01328_),
    .B(_01329_),
    .X(_01330_));
 sky130_fd_sc_hd__o2111a_1 _08713_ (.A1(_00955_),
    .A2(_00956_),
    .B1(_01322_),
    .C1(_01327_),
    .D1(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__buf_2 _08714_ (.A(net110),
    .X(_01332_));
 sky130_fd_sc_hd__and4_1 _08715_ (.A(_01332_),
    .B(_02334_),
    .C(_06611_),
    .D(_06602_),
    .X(_01333_));
 sky130_fd_sc_hd__a22oi_2 _08716_ (.A1(_06500_),
    .A2(_04778_),
    .B1(_04832_),
    .B2(_06501_),
    .Y(_01334_));
 sky130_fd_sc_hd__and4bb_1 _08717_ (.A_N(_01333_),
    .B_N(_01334_),
    .C(_06475_),
    .D(_00040_),
    .X(_01335_));
 sky130_fd_sc_hd__nor2_1 _08718_ (.A(_01333_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _08719_ (.A(_02528_),
    .B(_04585_),
    .Y(_01337_));
 sky130_fd_sc_hd__and4_1 _08720_ (.A(_06564_),
    .B(_02474_),
    .C(_00030_),
    .D(_00032_),
    .X(_01338_));
 sky130_fd_sc_hd__a22o_1 _08721_ (.A1(_02474_),
    .A2(_00030_),
    .B1(_00032_),
    .B2(_06564_),
    .X(_01339_));
 sky130_fd_sc_hd__and2b_1 _08722_ (.A_N(_01338_),
    .B(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__xnor2_1 _08723_ (.A(_01337_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__or2b_1 _08724_ (.A(_01336_),
    .B_N(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__a22o_1 _08725_ (.A1(_06515_),
    .A2(_04574_),
    .B1(_00030_),
    .B2(_06519_),
    .X(_01343_));
 sky130_fd_sc_hd__and4_1 _08726_ (.A(_06519_),
    .B(_06515_),
    .C(net6),
    .D(net7),
    .X(_01344_));
 sky130_fd_sc_hd__a31o_1 _08727_ (.A1(_02550_),
    .A2(_04531_),
    .A3(_01343_),
    .B1(_01344_),
    .X(_01345_));
 sky130_fd_sc_hd__xnor2_1 _08728_ (.A(_01336_),
    .B(_01341_),
    .Y(_01346_));
 sky130_fd_sc_hd__nand2_1 _08729_ (.A(_01345_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _08730_ (.A(_02712_),
    .B(_04445_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_2 _08731_ (.A(_06622_),
    .B(_04574_),
    .Y(_01349_));
 sky130_fd_sc_hd__nand2_2 _08732_ (.A(_00414_),
    .B(_04509_),
    .Y(_01350_));
 sky130_fd_sc_hd__a22o_1 _08733_ (.A1(_02647_),
    .A2(_00084_),
    .B1(_04574_),
    .B2(_02582_),
    .X(_01351_));
 sky130_fd_sc_hd__o21a_1 _08734_ (.A1(_01349_),
    .A2(_01350_),
    .B1(_01351_),
    .X(_01352_));
 sky130_fd_sc_hd__xnor2_1 _08735_ (.A(_01348_),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__and4_1 _08736_ (.A(_02582_),
    .B(_02647_),
    .C(_00082_),
    .D(_00084_),
    .X(_01354_));
 sky130_fd_sc_hd__a22oi_1 _08737_ (.A1(_06622_),
    .A2(_04434_),
    .B1(_00098_),
    .B2(_00414_),
    .Y(_01355_));
 sky130_fd_sc_hd__and4bb_1 _08738_ (.A_N(_01354_),
    .B_N(_01355_),
    .C(_06680_),
    .D(_00090_),
    .X(_01356_));
 sky130_fd_sc_hd__nor2_1 _08739_ (.A(_01354_),
    .B(_01356_),
    .Y(_01357_));
 sky130_fd_sc_hd__xnor2_1 _08740_ (.A(_01353_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__and4_1 _08741_ (.A(_06598_),
    .B(_06599_),
    .C(_04294_),
    .D(_00072_),
    .X(_01359_));
 sky130_fd_sc_hd__a22oi_1 _08742_ (.A1(_02797_),
    .A2(_00074_),
    .B1(_00090_),
    .B2(_02754_),
    .Y(_01360_));
 sky130_fd_sc_hd__and4bb_1 _08743_ (.A_N(_01359_),
    .B_N(_01360_),
    .C(_06608_),
    .D(_00301_),
    .X(_01361_));
 sky130_fd_sc_hd__o2bb2a_1 _08744_ (.A1_N(_02840_),
    .A2_N(_04251_),
    .B1(_01359_),
    .B2(_01360_),
    .X(_01362_));
 sky130_fd_sc_hd__nor2_1 _08745_ (.A(_01361_),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__xnor2_1 _08746_ (.A(_01358_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__a21o_2 _08747_ (.A1(_01342_),
    .A2(_01347_),
    .B1(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__and4_1 _08748_ (.A(_02582_),
    .B(_02647_),
    .C(_00089_),
    .D(_00082_),
    .X(_01366_));
 sky130_fd_sc_hd__a22oi_1 _08749_ (.A1(_06622_),
    .A2(_00072_),
    .B1(_00083_),
    .B2(_00414_),
    .Y(_01367_));
 sky130_fd_sc_hd__and4bb_1 _08750_ (.A_N(_01366_),
    .B_N(_01367_),
    .C(_06680_),
    .D(_00074_),
    .X(_01368_));
 sky130_fd_sc_hd__nor2_1 _08751_ (.A(_01366_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__o2bb2a_1 _08752_ (.A1_N(_06593_),
    .A2_N(_04369_),
    .B1(_01354_),
    .B2(_01355_),
    .X(_01370_));
 sky130_fd_sc_hd__nor2_1 _08753_ (.A(_01356_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__and2b_1 _08754_ (.A_N(_01369_),
    .B(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__xnor2_1 _08755_ (.A(_01371_),
    .B(_01369_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _08756_ (.A(_06608_),
    .B(_00272_),
    .Y(_01374_));
 sky130_fd_sc_hd__and4_1 _08757_ (.A(_06606_),
    .B(_06601_),
    .C(_04240_),
    .D(_00074_),
    .X(_01375_));
 sky130_fd_sc_hd__a22oi_2 _08758_ (.A1(_00878_),
    .A2(_00301_),
    .B1(_00259_),
    .B2(_00877_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _08759_ (.A(_01375_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__xnor2_2 _08760_ (.A(_01374_),
    .B(_01377_),
    .Y(_01378_));
 sky130_fd_sc_hd__and2_1 _08761_ (.A(_01373_),
    .B(_01378_),
    .X(_01379_));
 sky130_fd_sc_hd__nand3_2 _08762_ (.A(_01342_),
    .B(_01347_),
    .C(_01364_),
    .Y(_01380_));
 sky130_fd_sc_hd__o211ai_4 _08763_ (.A1(_01372_),
    .A2(_01379_),
    .B1(_01380_),
    .C1(_01365_),
    .Y(_01381_));
 sky130_fd_sc_hd__o21ba_1 _08764_ (.A1(_01374_),
    .A2(_01376_),
    .B1_N(_01375_),
    .X(_01382_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_03002_),
    .B(_06443_),
    .Y(_01383_));
 sky130_fd_sc_hd__and4_1 _08766_ (.A(net120),
    .B(net44),
    .C(_04100_),
    .D(_04165_),
    .X(_01384_));
 sky130_fd_sc_hd__a22o_1 _08767_ (.A1(_00029_),
    .A2(_04100_),
    .B1(_00271_),
    .B2(net120),
    .X(_01385_));
 sky130_fd_sc_hd__and2b_1 _08768_ (.A_N(_01384_),
    .B(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__xnor2_2 _08769_ (.A(_01383_),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__or2b_1 _08770_ (.A(_01382_),
    .B_N(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__a22o_1 _08771_ (.A1(_02948_),
    .A2(_06430_),
    .B1(_06431_),
    .B2(_00028_),
    .X(_01389_));
 sky130_fd_sc_hd__and4_1 _08772_ (.A(_00028_),
    .B(_00029_),
    .C(_06430_),
    .D(_06431_),
    .X(_01390_));
 sky130_fd_sc_hd__a31o_2 _08773_ (.A1(_03024_),
    .A2(_03982_),
    .A3(_01389_),
    .B1(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__xnor2_1 _08774_ (.A(_01382_),
    .B(_01387_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _08775_ (.A(_01391_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__a31o_2 _08776_ (.A1(_03024_),
    .A2(_04057_),
    .A3(_01385_),
    .B1(_01384_),
    .X(_01394_));
 sky130_fd_sc_hd__nor2_1 _08777_ (.A(_01359_),
    .B(_01361_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_03002_),
    .B(_00303_),
    .Y(_01396_));
 sky130_fd_sc_hd__and4_1 _08779_ (.A(net120),
    .B(net44),
    .C(_00271_),
    .D(_04229_),
    .X(_01397_));
 sky130_fd_sc_hd__a22o_1 _08780_ (.A1(_00029_),
    .A2(_00271_),
    .B1(_04229_),
    .B2(_00028_),
    .X(_01398_));
 sky130_fd_sc_hd__and2b_1 _08781_ (.A_N(_01397_),
    .B(_01398_),
    .X(_01399_));
 sky130_fd_sc_hd__xnor2_2 _08782_ (.A(_01396_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__xnor2_1 _08783_ (.A(_01395_),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__xnor2_2 _08784_ (.A(_01394_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__a21oi_4 _08785_ (.A1(_01388_),
    .A2(_01393_),
    .B1(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__and3_1 _08786_ (.A(_01402_),
    .B(_01388_),
    .C(_01393_),
    .X(_01404_));
 sky130_fd_sc_hd__and4_1 _08787_ (.A(_00921_),
    .B(_01206_),
    .C(_03960_),
    .D(_06446_),
    .X(_01405_));
 sky130_fd_sc_hd__a22oi_1 _08788_ (.A1(_03110_),
    .A2(_06437_),
    .B1(_04046_),
    .B2(_03067_),
    .Y(_01406_));
 sky130_fd_sc_hd__and4bb_1 _08789_ (.A_N(_01405_),
    .B_N(_01406_),
    .C(_03174_),
    .D(_03884_),
    .X(_01407_));
 sky130_fd_sc_hd__nand4_4 _08790_ (.A(_03067_),
    .B(_03110_),
    .C(_03895_),
    .D(_03993_),
    .Y(_01408_));
 sky130_fd_sc_hd__o2bb2a_1 _08791_ (.A1_N(_03174_),
    .A2_N(_03895_),
    .B1(_01405_),
    .B2(_01406_),
    .X(_01409_));
 sky130_fd_sc_hd__nor3_1 _08792_ (.A(_01407_),
    .B(_01408_),
    .C(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__o21a_1 _08793_ (.A1(_01407_),
    .A2(_01409_),
    .B1(_01408_),
    .X(_01411_));
 sky130_fd_sc_hd__or2_1 _08794_ (.A(_01410_),
    .B(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__nor3_4 _08795_ (.A(_01403_),
    .B(_01404_),
    .C(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__o21a_1 _08796_ (.A1(_01403_),
    .A2(_01404_),
    .B1(_01412_),
    .X(_01414_));
 sky130_fd_sc_hd__a211oi_4 _08797_ (.A1(_01365_),
    .A2(_01381_),
    .B1(_01413_),
    .C1(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__and4_1 _08798_ (.A(_02754_),
    .B(_02797_),
    .C(_00287_),
    .D(_00267_),
    .X(_01416_));
 sky130_fd_sc_hd__a22oi_1 _08799_ (.A1(_06630_),
    .A2(_04176_),
    .B1(_04240_),
    .B2(_06631_),
    .Y(_01417_));
 sky130_fd_sc_hd__and4bb_1 _08800_ (.A_N(_01416_),
    .B_N(_01417_),
    .C(_06608_),
    .D(_00303_),
    .X(_01418_));
 sky130_fd_sc_hd__nor2_2 _08801_ (.A(_01416_),
    .B(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__nand2_2 _08802_ (.A(_00444_),
    .B(_06437_),
    .Y(_01420_));
 sky130_fd_sc_hd__and2b_1 _08803_ (.A_N(_01390_),
    .B(_01389_),
    .X(_01421_));
 sky130_fd_sc_hd__xnor2_4 _08804_ (.A(_01420_),
    .B(_01421_),
    .Y(_01422_));
 sky130_fd_sc_hd__or2b_1 _08805_ (.A(_01419_),
    .B_N(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__and4_1 _08806_ (.A(_00049_),
    .B(_00062_),
    .C(_06436_),
    .D(_04035_),
    .X(_01424_));
 sky130_fd_sc_hd__a22oi_1 _08807_ (.A1(_02959_),
    .A2(_03960_),
    .B1(_06443_),
    .B2(_02905_),
    .Y(_01425_));
 sky130_fd_sc_hd__and4bb_1 _08808_ (.A_N(_01424_),
    .B_N(_01425_),
    .C(_00444_),
    .D(_03873_),
    .X(_01426_));
 sky130_fd_sc_hd__or2_2 _08809_ (.A(_01424_),
    .B(_01426_),
    .X(_01427_));
 sky130_fd_sc_hd__xnor2_1 _08810_ (.A(_01419_),
    .B(_01422_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(_01427_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__xnor2_1 _08812_ (.A(_01391_),
    .B(_01392_),
    .Y(_01430_));
 sky130_fd_sc_hd__a21o_1 _08813_ (.A1(_01423_),
    .A2(_01429_),
    .B1(_01430_),
    .X(_01431_));
 sky130_fd_sc_hd__nand3_1 _08814_ (.A(_01430_),
    .B(_01423_),
    .C(_01429_),
    .Y(_01432_));
 sky130_fd_sc_hd__a22o_1 _08815_ (.A1(_03110_),
    .A2(_03906_),
    .B1(_03993_),
    .B2(_03067_),
    .X(_01433_));
 sky130_fd_sc_hd__nand4_2 _08816_ (.A(_01408_),
    .B(_01431_),
    .C(_01432_),
    .D(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__o211a_1 _08817_ (.A1(_01413_),
    .A2(_01414_),
    .B1(_01365_),
    .C1(_01381_),
    .X(_01435_));
 sky130_fd_sc_hd__a211oi_2 _08818_ (.A1(_01431_),
    .A2(_01434_),
    .B1(_01435_),
    .C1(_01415_),
    .Y(_01436_));
 sky130_fd_sc_hd__o21ai_2 _08819_ (.A1(_01415_),
    .A2(_01436_),
    .B1(_01410_),
    .Y(_01437_));
 sky130_fd_sc_hd__and4_1 _08820_ (.A(_02096_),
    .B(_02194_),
    .C(net14),
    .D(net15),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(net111),
    .B(_06581_),
    .Y(_01439_));
 sky130_fd_sc_hd__a22oi_2 _08822_ (.A1(_00150_),
    .A2(net14),
    .B1(_05176_),
    .B2(_06494_),
    .Y(_01440_));
 sky130_fd_sc_hd__or3_1 _08823_ (.A(_01438_),
    .B(_01439_),
    .C(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__nand2_1 _08824_ (.A(_06460_),
    .B(net133),
    .Y(_01442_));
 sky130_fd_sc_hd__a22oi_2 _08825_ (.A1(_06495_),
    .A2(_06581_),
    .B1(_05101_),
    .B2(_02107_),
    .Y(_01443_));
 sky130_fd_sc_hd__and4_1 _08826_ (.A(_02096_),
    .B(_02194_),
    .C(net13),
    .D(net14),
    .X(_01444_));
 sky130_fd_sc_hd__o21bai_1 _08827_ (.A1(_01442_),
    .A2(_01443_),
    .B1_N(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__o21ai_1 _08828_ (.A1(_01438_),
    .A2(_01440_),
    .B1(_01439_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand3_1 _08829_ (.A(_01441_),
    .B(_01445_),
    .C(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__a21o_1 _08830_ (.A1(_01441_),
    .A2(_01446_),
    .B1(_01445_),
    .X(_01448_));
 sky130_fd_sc_hd__nand2_1 _08831_ (.A(_06544_),
    .B(_06603_),
    .Y(_01449_));
 sky130_fd_sc_hd__a22oi_2 _08832_ (.A1(_06548_),
    .A2(_04896_),
    .B1(_04961_),
    .B2(_02291_),
    .Y(_01450_));
 sky130_fd_sc_hd__and4_1 _08833_ (.A(_01332_),
    .B(_02334_),
    .C(_06604_),
    .D(_06580_),
    .X(_01451_));
 sky130_fd_sc_hd__nor2_1 _08834_ (.A(_01450_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__xnor2_1 _08835_ (.A(_01449_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand3_1 _08836_ (.A(_01447_),
    .B(_01448_),
    .C(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__or3_1 _08837_ (.A(_01444_),
    .B(_01442_),
    .C(_01443_),
    .X(_01455_));
 sky130_fd_sc_hd__o21ai_1 _08838_ (.A1(_01444_),
    .A2(_01443_),
    .B1(_01442_),
    .Y(_01456_));
 sky130_fd_sc_hd__and2_1 _08839_ (.A(_06460_),
    .B(_06604_),
    .X(_01457_));
 sky130_fd_sc_hd__a22o_1 _08840_ (.A1(_06463_),
    .A2(net133),
    .B1(_06581_),
    .B2(_02107_),
    .X(_01458_));
 sky130_fd_sc_hd__nand4_1 _08841_ (.A(_06534_),
    .B(_06491_),
    .C(_06580_),
    .D(_06581_),
    .Y(_01459_));
 sky130_fd_sc_hd__a21bo_1 _08842_ (.A1(_01457_),
    .A2(_01458_),
    .B1_N(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__a21o_1 _08843_ (.A1(_01455_),
    .A2(_01456_),
    .B1(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(_06544_),
    .B(_04778_),
    .Y(_01462_));
 sky130_fd_sc_hd__a22oi_1 _08845_ (.A1(_06548_),
    .A2(_04832_),
    .B1(_04896_),
    .B2(_02291_),
    .Y(_01463_));
 sky130_fd_sc_hd__and4_1 _08846_ (.A(_01332_),
    .B(_02334_),
    .C(_06602_),
    .D(_06604_),
    .X(_01464_));
 sky130_fd_sc_hd__nor2_1 _08847_ (.A(_01463_),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__xnor2_1 _08848_ (.A(_01462_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand3_1 _08849_ (.A(_01455_),
    .B(_01460_),
    .C(_01456_),
    .Y(_01467_));
 sky130_fd_sc_hd__a21bo_1 _08850_ (.A1(_01461_),
    .A2(_01466_),
    .B1_N(_01467_),
    .X(_01468_));
 sky130_fd_sc_hd__a21o_1 _08851_ (.A1(_01447_),
    .A2(_01448_),
    .B1(_01453_),
    .X(_01469_));
 sky130_fd_sc_hd__nand3_2 _08852_ (.A(_01454_),
    .B(_01468_),
    .C(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hd__a21o_1 _08853_ (.A1(_01454_),
    .A2(_01469_),
    .B1(_01468_),
    .X(_01471_));
 sky130_fd_sc_hd__a31o_1 _08854_ (.A1(_02539_),
    .A2(_04596_),
    .A3(_01339_),
    .B1(_01338_),
    .X(_01472_));
 sky130_fd_sc_hd__o21ba_1 _08855_ (.A1(_01462_),
    .A2(_01463_),
    .B1_N(_01464_),
    .X(_01473_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_06663_),
    .B(_00048_),
    .Y(_01474_));
 sky130_fd_sc_hd__and4_1 _08857_ (.A(net107),
    .B(net66),
    .C(net8),
    .D(_04767_),
    .X(_01475_));
 sky130_fd_sc_hd__a22o_1 _08858_ (.A1(_06515_),
    .A2(_00032_),
    .B1(_04767_),
    .B2(net107),
    .X(_01476_));
 sky130_fd_sc_hd__and2b_1 _08859_ (.A_N(_01475_),
    .B(_01476_),
    .X(_01477_));
 sky130_fd_sc_hd__xnor2_2 _08860_ (.A(_01474_),
    .B(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__xnor2_1 _08861_ (.A(_01473_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__xor2_1 _08862_ (.A(_01472_),
    .B(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__nand3_1 _08863_ (.A(_01470_),
    .B(_01471_),
    .C(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__or3_1 _08864_ (.A(_01283_),
    .B(_01281_),
    .C(_01282_),
    .X(_01482_));
 sky130_fd_sc_hd__o21bai_1 _08865_ (.A1(_01439_),
    .A2(_01440_),
    .B1_N(_01438_),
    .Y(_01483_));
 sky130_fd_sc_hd__o21ai_1 _08866_ (.A1(_01283_),
    .A2(_01282_),
    .B1(_01281_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand3_1 _08867_ (.A(_01482_),
    .B(_01483_),
    .C(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__a21o_1 _08868_ (.A1(_01482_),
    .A2(_01484_),
    .B1(_01483_),
    .X(_01486_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_06475_),
    .B(_04907_),
    .Y(_01487_));
 sky130_fd_sc_hd__a22oi_1 _08870_ (.A1(_06500_),
    .A2(_06580_),
    .B1(_05025_),
    .B2(_06501_),
    .Y(_01488_));
 sky130_fd_sc_hd__and4_1 _08871_ (.A(_06503_),
    .B(_06504_),
    .C(_06580_),
    .D(_06581_),
    .X(_01489_));
 sky130_fd_sc_hd__nor2_1 _08872_ (.A(_01488_),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__xnor2_1 _08873_ (.A(_01487_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand3_1 _08874_ (.A(_01485_),
    .B(_01486_),
    .C(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__a21bo_1 _08875_ (.A1(_01448_),
    .A2(_01453_),
    .B1_N(_01447_),
    .X(_01493_));
 sky130_fd_sc_hd__a21o_1 _08876_ (.A1(_01485_),
    .A2(_01486_),
    .B1(_01491_),
    .X(_01494_));
 sky130_fd_sc_hd__nand3_2 _08877_ (.A(_01492_),
    .B(_01493_),
    .C(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__a21o_1 _08878_ (.A1(_01492_),
    .A2(_01494_),
    .B1(_01493_),
    .X(_01496_));
 sky130_fd_sc_hd__a31o_1 _08879_ (.A1(_02539_),
    .A2(_04660_),
    .A3(_01476_),
    .B1(_01475_),
    .X(_01497_));
 sky130_fd_sc_hd__o21ba_1 _08880_ (.A1(_01449_),
    .A2(_01450_),
    .B1_N(_01451_),
    .X(_01498_));
 sky130_fd_sc_hd__and4_1 _08881_ (.A(_06519_),
    .B(_06515_),
    .C(_04767_),
    .D(net10),
    .X(_01499_));
 sky130_fd_sc_hd__a22oi_1 _08882_ (.A1(_06513_),
    .A2(_06611_),
    .B1(_04832_),
    .B2(_02420_),
    .Y(_01500_));
 sky130_fd_sc_hd__and4bb_1 _08883_ (.A_N(_01499_),
    .B_N(_01500_),
    .C(_06663_),
    .D(_00033_),
    .X(_01501_));
 sky130_fd_sc_hd__o2bb2a_1 _08884_ (.A1_N(_06663_),
    .A2_N(_00033_),
    .B1(_01499_),
    .B2(_01500_),
    .X(_01502_));
 sky130_fd_sc_hd__nor2_1 _08885_ (.A(_01501_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(_01498_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__xor2_1 _08887_ (.A(_01497_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__a21oi_1 _08888_ (.A1(_01495_),
    .A2(_01496_),
    .B1(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__and3_1 _08889_ (.A(_01495_),
    .B(_01496_),
    .C(_01505_),
    .X(_01507_));
 sky130_fd_sc_hd__a211oi_2 _08890_ (.A1(_01470_),
    .A2(_01481_),
    .B1(_01506_),
    .C1(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__o211a_1 _08891_ (.A1(_01507_),
    .A2(_01506_),
    .B1(_01481_),
    .C1(_01470_),
    .X(_01509_));
 sky130_fd_sc_hd__and2b_1 _08892_ (.A_N(_01357_),
    .B(_01353_),
    .X(_01510_));
 sky130_fd_sc_hd__and2_1 _08893_ (.A(_01358_),
    .B(_01363_),
    .X(_01511_));
 sky130_fd_sc_hd__or2b_1 _08894_ (.A(_01473_),
    .B_N(_01478_),
    .X(_01512_));
 sky130_fd_sc_hd__nand2_1 _08895_ (.A(_01472_),
    .B(_01479_),
    .Y(_01513_));
 sky130_fd_sc_hd__and4_1 _08896_ (.A(_06578_),
    .B(_02647_),
    .C(_04574_),
    .D(_00030_),
    .X(_01514_));
 sky130_fd_sc_hd__a22oi_1 _08897_ (.A1(_06622_),
    .A2(_00035_),
    .B1(_04638_),
    .B2(_00414_),
    .Y(_01515_));
 sky130_fd_sc_hd__and4bb_1 _08898_ (.A_N(_01514_),
    .B_N(_01515_),
    .C(_06680_),
    .D(_00085_),
    .X(_01516_));
 sky130_fd_sc_hd__o2bb2a_1 _08899_ (.A1_N(_06593_),
    .A2_N(_04520_),
    .B1(_01514_),
    .B2(_01515_),
    .X(_01517_));
 sky130_fd_sc_hd__nor2_1 _08900_ (.A(_01516_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _08901_ (.A(_01349_),
    .B(_01350_),
    .Y(_01519_));
 sky130_fd_sc_hd__a31o_1 _08902_ (.A1(_06620_),
    .A2(_04456_),
    .A3(_01351_),
    .B1(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__xor2_1 _08903_ (.A(_01518_),
    .B(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__and4_1 _08904_ (.A(_02754_),
    .B(_02797_),
    .C(_04358_),
    .D(_00083_),
    .X(_01522_));
 sky130_fd_sc_hd__a22oi_1 _08905_ (.A1(_06630_),
    .A2(_00090_),
    .B1(_00093_),
    .B2(_06631_),
    .Y(_01523_));
 sky130_fd_sc_hd__and4bb_1 _08906_ (.A_N(_01522_),
    .B_N(_01523_),
    .C(_06608_),
    .D(_00259_),
    .X(_01524_));
 sky130_fd_sc_hd__o2bb2a_1 _08907_ (.A1_N(_06610_),
    .A2_N(_04316_),
    .B1(_01522_),
    .B2(_01523_),
    .X(_01525_));
 sky130_fd_sc_hd__nor2_1 _08908_ (.A(_01524_),
    .B(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__xnor2_1 _08909_ (.A(_01521_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__a21o_1 _08910_ (.A1(_01512_),
    .A2(_01513_),
    .B1(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__nand3_1 _08911_ (.A(_01512_),
    .B(_01513_),
    .C(_01527_),
    .Y(_01529_));
 sky130_fd_sc_hd__o211ai_2 _08912_ (.A1(_01510_),
    .A2(_01511_),
    .B1(_01528_),
    .C1(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__a211o_1 _08913_ (.A1(_01528_),
    .A2(_01529_),
    .B1(_01510_),
    .C1(_01511_),
    .X(_01531_));
 sky130_fd_sc_hd__and4bb_1 _08914_ (.A_N(_01508_),
    .B_N(_01509_),
    .C(_01530_),
    .D(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__nand3_1 _08915_ (.A(_01495_),
    .B(_01496_),
    .C(_01505_),
    .Y(_01533_));
 sky130_fd_sc_hd__nand3_1 _08916_ (.A(_01288_),
    .B(_01285_),
    .C(_01287_),
    .Y(_01534_));
 sky130_fd_sc_hd__a21bo_1 _08917_ (.A1(_01486_),
    .A2(_01491_),
    .B1_N(_01485_),
    .X(_01535_));
 sky130_fd_sc_hd__a21o_1 _08918_ (.A1(_01288_),
    .A2(_01285_),
    .B1(_01287_),
    .X(_01536_));
 sky130_fd_sc_hd__nand3_2 _08919_ (.A(_01534_),
    .B(_01535_),
    .C(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__a21o_1 _08920_ (.A1(_01534_),
    .A2(_01536_),
    .B1(_01535_),
    .X(_01538_));
 sky130_fd_sc_hd__nor2_1 _08921_ (.A(_01499_),
    .B(_01501_),
    .Y(_01539_));
 sky130_fd_sc_hd__o21ba_1 _08922_ (.A1(_01487_),
    .A2(_01488_),
    .B1_N(_01489_),
    .X(_01540_));
 sky130_fd_sc_hd__nand2_1 _08923_ (.A(_06560_),
    .B(_04789_),
    .Y(_01541_));
 sky130_fd_sc_hd__xnor2_1 _08924_ (.A(_01541_),
    .B(_01217_),
    .Y(_01542_));
 sky130_fd_sc_hd__xnor2_1 _08925_ (.A(_01540_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__xnor2_1 _08926_ (.A(_01539_),
    .B(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__a21oi_1 _08927_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__and3_1 _08928_ (.A(_01537_),
    .B(_01538_),
    .C(_01544_),
    .X(_01546_));
 sky130_fd_sc_hd__a211oi_2 _08929_ (.A1(_01495_),
    .A2(_01533_),
    .B1(_01545_),
    .C1(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__o211a_1 _08930_ (.A1(_01546_),
    .A2(_01545_),
    .B1(_01533_),
    .C1(_01495_),
    .X(_01548_));
 sky130_fd_sc_hd__and2_1 _08931_ (.A(_01518_),
    .B(_01520_),
    .X(_01549_));
 sky130_fd_sc_hd__and2_1 _08932_ (.A(_01521_),
    .B(_01526_),
    .X(_01550_));
 sky130_fd_sc_hd__or3_1 _08933_ (.A(_01501_),
    .B(_01498_),
    .C(_01502_),
    .X(_01551_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(_01497_),
    .B(_01504_),
    .Y(_01552_));
 sky130_fd_sc_hd__o2bb2a_1 _08935_ (.A1_N(_06620_),
    .A2_N(_00036_),
    .B1(_01229_),
    .B2(_01230_),
    .X(_01553_));
 sky130_fd_sc_hd__nor2_1 _08936_ (.A(_01231_),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__nor2_1 _08937_ (.A(_01514_),
    .B(_01516_),
    .Y(_01555_));
 sky130_fd_sc_hd__xnor2_1 _08938_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__o2bb2a_1 _08939_ (.A1_N(_02851_),
    .A2_N(_04380_),
    .B1(_01246_),
    .B2(_01247_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _08940_ (.A(_01248_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__xnor2_1 _08941_ (.A(_01556_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__a21o_1 _08942_ (.A1(_01551_),
    .A2(_01552_),
    .B1(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__nand3_1 _08943_ (.A(_01551_),
    .B(_01552_),
    .C(_01559_),
    .Y(_01561_));
 sky130_fd_sc_hd__o211ai_2 _08944_ (.A1(_01549_),
    .A2(_01550_),
    .B1(_01560_),
    .C1(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__a211o_1 _08945_ (.A1(_01560_),
    .A2(_01561_),
    .B1(_01549_),
    .C1(_01550_),
    .X(_01563_));
 sky130_fd_sc_hd__a2bb2o_1 _08946_ (.A1_N(_01547_),
    .A2_N(_01548_),
    .B1(_01562_),
    .B2(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__or4bb_1 _08947_ (.A(_01547_),
    .B(_01548_),
    .C_N(_01562_),
    .D_N(_01563_),
    .X(_01565_));
 sky130_fd_sc_hd__o211a_1 _08948_ (.A1(_01508_),
    .A2(_01532_),
    .B1(_01564_),
    .C1(_01565_),
    .X(_01566_));
 sky130_fd_sc_hd__a211oi_1 _08949_ (.A1(_01565_),
    .A2(_01564_),
    .B1(_01532_),
    .C1(_01508_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2b_1 _08950_ (.A(_01395_),
    .B_N(_01400_),
    .X(_01568_));
 sky130_fd_sc_hd__nand2_1 _08951_ (.A(_01394_),
    .B(_01401_),
    .Y(_01569_));
 sky130_fd_sc_hd__a31o_1 _08952_ (.A1(_03024_),
    .A2(_04122_),
    .A3(_01398_),
    .B1(_01397_),
    .X(_01570_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_01522_),
    .B(_01524_),
    .Y(_01571_));
 sky130_fd_sc_hd__o2bb2a_1 _08954_ (.A1_N(_00058_),
    .A2_N(_00272_),
    .B1(_01253_),
    .B2(_01254_),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_1 _08955_ (.A(_01255_),
    .B(_01572_),
    .Y(_01573_));
 sky130_fd_sc_hd__xnor2_1 _08956_ (.A(_01571_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__xnor2_1 _08957_ (.A(_01570_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__a21o_1 _08958_ (.A1(_01568_),
    .A2(_01569_),
    .B1(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__nand3_1 _08959_ (.A(_01575_),
    .B(_01568_),
    .C(_01569_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_03239_),
    .B(_03906_),
    .Y(_01578_));
 sky130_fd_sc_hd__a22oi_1 _08961_ (.A1(_03174_),
    .A2(_03971_),
    .B1(_01205_),
    .B2(_01207_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _08962_ (.A(_01208_),
    .B(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_01405_),
    .B(_01407_),
    .Y(_01581_));
 sky130_fd_sc_hd__xnor2_1 _08964_ (.A(_01580_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__xnor2_1 _08965_ (.A(_01578_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__a21oi_1 _08966_ (.A1(_01576_),
    .A2(_01577_),
    .B1(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__and3_1 _08967_ (.A(_01576_),
    .B(_01577_),
    .C(_01583_),
    .X(_01585_));
 sky130_fd_sc_hd__a211o_1 _08968_ (.A1(_01528_),
    .A2(_01530_),
    .B1(_01584_),
    .C1(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__o211ai_2 _08969_ (.A1(_01585_),
    .A2(_01584_),
    .B1(_01530_),
    .C1(_01528_),
    .Y(_01587_));
 sky130_fd_sc_hd__o211ai_2 _08970_ (.A1(_01403_),
    .A2(_01413_),
    .B1(_01586_),
    .C1(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__a211o_1 _08971_ (.A1(_01586_),
    .A2(_01587_),
    .B1(_01403_),
    .C1(_01413_),
    .X(_01589_));
 sky130_fd_sc_hd__and4bb_1 _08972_ (.A_N(_01566_),
    .B_N(_01567_),
    .C(_01588_),
    .D(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__a2bb2oi_1 _08973_ (.A1_N(_01566_),
    .A2_N(_01567_),
    .B1(_01588_),
    .B2(_01589_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand3_1 _08974_ (.A(_01457_),
    .B(_01459_),
    .C(_01458_),
    .Y(_01592_));
 sky130_fd_sc_hd__a21o_1 _08975_ (.A1(_01459_),
    .A2(_01458_),
    .B1(_01457_),
    .X(_01593_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(_06488_),
    .B(_04832_),
    .Y(_01594_));
 sky130_fd_sc_hd__a22oi_2 _08977_ (.A1(_06491_),
    .A2(_06604_),
    .B1(_06580_),
    .B2(_06492_),
    .Y(_01595_));
 sky130_fd_sc_hd__and4_1 _08978_ (.A(_06494_),
    .B(_06495_),
    .C(net11),
    .D(net133),
    .X(_01596_));
 sky130_fd_sc_hd__o21bai_1 _08979_ (.A1(_01594_),
    .A2(_01595_),
    .B1_N(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21o_1 _08980_ (.A1(_01592_),
    .A2(_01593_),
    .B1(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__o2bb2a_1 _08981_ (.A1_N(_02377_),
    .A2_N(_04714_),
    .B1(_01333_),
    .B2(_01334_),
    .X(_01599_));
 sky130_fd_sc_hd__nor2_1 _08982_ (.A(_01335_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__nand3_1 _08983_ (.A(_01597_),
    .B(_01592_),
    .C(_01593_),
    .Y(_01601_));
 sky130_fd_sc_hd__a21bo_1 _08984_ (.A1(_01598_),
    .A2(_01600_),
    .B1_N(_01601_),
    .X(_01602_));
 sky130_fd_sc_hd__nand3_1 _08985_ (.A(_01467_),
    .B(_01461_),
    .C(_01466_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21o_1 _08986_ (.A1(_01467_),
    .A2(_01461_),
    .B1(_01466_),
    .X(_01604_));
 sky130_fd_sc_hd__nand3_2 _08987_ (.A(_01602_),
    .B(_01603_),
    .C(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__a21o_1 _08988_ (.A1(_01603_),
    .A2(_01604_),
    .B1(_01602_),
    .X(_01606_));
 sky130_fd_sc_hd__xor2_1 _08989_ (.A(_01345_),
    .B(_01346_),
    .X(_01607_));
 sky130_fd_sc_hd__nand3_1 _08990_ (.A(_01605_),
    .B(_01606_),
    .C(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__and3_1 _08991_ (.A(_01470_),
    .B(_01471_),
    .C(_01480_),
    .X(_01609_));
 sky130_fd_sc_hd__a21oi_1 _08992_ (.A1(_01470_),
    .A2(_01471_),
    .B1(_01480_),
    .Y(_01610_));
 sky130_fd_sc_hd__a211oi_2 _08993_ (.A1(_01605_),
    .A2(_01608_),
    .B1(_01609_),
    .C1(_01610_),
    .Y(_01611_));
 sky130_fd_sc_hd__o211a_1 _08994_ (.A1(_01372_),
    .A2(_01379_),
    .B1(_01380_),
    .C1(_01365_),
    .X(_01612_));
 sky130_fd_sc_hd__o211a_1 _08995_ (.A1(_01609_),
    .A2(_01610_),
    .B1(_01605_),
    .C1(_01608_),
    .X(_01613_));
 sky130_fd_sc_hd__a211o_1 _08996_ (.A1(_01365_),
    .A2(_01380_),
    .B1(_01379_),
    .C1(_01372_),
    .X(_01614_));
 sky130_fd_sc_hd__nor4b_1 _08997_ (.A(_01612_),
    .B(_01611_),
    .C(_01613_),
    .D_N(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__or4bb_1 _08998_ (.A(_01508_),
    .B(_01509_),
    .C_N(_01530_),
    .D_N(_01531_),
    .X(_01616_));
 sky130_fd_sc_hd__a2bb2o_1 _08999_ (.A1_N(_01508_),
    .A2_N(_01509_),
    .B1(_01530_),
    .B2(_01531_),
    .X(_01617_));
 sky130_fd_sc_hd__o211ai_2 _09000_ (.A1(_01611_),
    .A2(_01615_),
    .B1(_01616_),
    .C1(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__a211o_1 _09001_ (.A1(_01616_),
    .A2(_01617_),
    .B1(_01611_),
    .C1(_01615_),
    .X(_01619_));
 sky130_fd_sc_hd__o211ai_1 _09002_ (.A1(_01415_),
    .A2(_01435_),
    .B1(_01434_),
    .C1(_01431_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand4b_1 _09003_ (.A_N(_01436_),
    .B(_01618_),
    .C(_01619_),
    .D(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__o211ai_1 _09004_ (.A1(_01590_),
    .A2(_01591_),
    .B1(_01618_),
    .C1(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__or3_1 _09005_ (.A(_01410_),
    .B(_01415_),
    .C(_01436_),
    .X(_01623_));
 sky130_fd_sc_hd__and2_1 _09006_ (.A(_01437_),
    .B(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__a211o_1 _09007_ (.A1(_01618_),
    .A2(_01621_),
    .B1(_01590_),
    .C1(_01591_),
    .X(_01625_));
 sky130_fd_sc_hd__a21boi_1 _09008_ (.A1(_01622_),
    .A2(_01624_),
    .B1_N(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__and4bb_1 _09009_ (.A_N(_01547_),
    .B_N(_01548_),
    .C(_01562_),
    .D(_01563_),
    .X(_01627_));
 sky130_fd_sc_hd__nand3_1 _09010_ (.A(_01537_),
    .B(_01538_),
    .C(_01544_),
    .Y(_01628_));
 sky130_fd_sc_hd__a21oi_2 _09011_ (.A1(_01291_),
    .A2(_01292_),
    .B1(_01294_),
    .Y(_01629_));
 sky130_fd_sc_hd__and3_1 _09012_ (.A(_01291_),
    .B(_01292_),
    .C(_01294_),
    .X(_01630_));
 sky130_fd_sc_hd__a211oi_4 _09013_ (.A1(_01537_),
    .A2(_01628_),
    .B1(_01629_),
    .C1(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__o211a_1 _09014_ (.A1(_01630_),
    .A2(_01629_),
    .B1(_01628_),
    .C1(_01537_),
    .X(_01632_));
 sky130_fd_sc_hd__and2b_1 _09015_ (.A_N(_01555_),
    .B(_01554_),
    .X(_01633_));
 sky130_fd_sc_hd__and2_1 _09016_ (.A(_01556_),
    .B(_01558_),
    .X(_01634_));
 sky130_fd_sc_hd__or2b_1 _09017_ (.A(_01540_),
    .B_N(_01542_),
    .X(_01635_));
 sky130_fd_sc_hd__or2b_1 _09018_ (.A(_01539_),
    .B_N(_01543_),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_1 _09019_ (.A(_01237_),
    .B(_01239_),
    .Y(_01637_));
 sky130_fd_sc_hd__a21o_1 _09020_ (.A1(_01635_),
    .A2(_01636_),
    .B1(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__nand3_1 _09021_ (.A(_01635_),
    .B(_01636_),
    .C(_01637_),
    .Y(_01639_));
 sky130_fd_sc_hd__o211ai_2 _09022_ (.A1(_01633_),
    .A2(_01634_),
    .B1(_01638_),
    .C1(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__a211o_1 _09023_ (.A1(_01638_),
    .A2(_01639_),
    .B1(_01633_),
    .C1(_01634_),
    .X(_01641_));
 sky130_fd_sc_hd__a2bb2o_1 _09024_ (.A1_N(_01631_),
    .A2_N(_01632_),
    .B1(_01640_),
    .B2(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__or4bb_1 _09025_ (.A(_01631_),
    .B(_01632_),
    .C_N(_01640_),
    .D_N(_01641_),
    .X(_01643_));
 sky130_fd_sc_hd__o211a_1 _09026_ (.A1(_01547_),
    .A2(_01627_),
    .B1(_01642_),
    .C1(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__a211oi_1 _09027_ (.A1(_01643_),
    .A2(_01642_),
    .B1(_01627_),
    .C1(_01547_),
    .Y(_01645_));
 sky130_fd_sc_hd__inv_2 _09028_ (.A(_01576_),
    .Y(_01646_));
 sky130_fd_sc_hd__or3_1 _09029_ (.A(_01255_),
    .B(_01571_),
    .C(_01572_),
    .X(_01647_));
 sky130_fd_sc_hd__nand2_1 _09030_ (.A(_01570_),
    .B(_01574_),
    .Y(_01648_));
 sky130_fd_sc_hd__xnor2_1 _09031_ (.A(_01256_),
    .B(_01257_),
    .Y(_01649_));
 sky130_fd_sc_hd__a21o_1 _09032_ (.A1(_01647_),
    .A2(_01648_),
    .B1(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__nand3_1 _09033_ (.A(_01649_),
    .B(_01647_),
    .C(_01648_),
    .Y(_01651_));
 sky130_fd_sc_hd__a22oi_2 _09034_ (.A1(_03293_),
    .A2(_03895_),
    .B1(_03982_),
    .B2(_03239_),
    .Y(_01652_));
 sky130_fd_sc_hd__or2_1 _09035_ (.A(_01203_),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__nor2_1 _09036_ (.A(_01204_),
    .B(_01208_),
    .Y(_01654_));
 sky130_fd_sc_hd__xnor2_2 _09037_ (.A(_01210_),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_1 _09038_ (.A(_01653_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__a21oi_1 _09039_ (.A1(_01650_),
    .A2(_01651_),
    .B1(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__and3_1 _09040_ (.A(_01650_),
    .B(_01651_),
    .C(_01656_),
    .X(_01658_));
 sky130_fd_sc_hd__a211o_1 _09041_ (.A1(_01560_),
    .A2(_01562_),
    .B1(_01657_),
    .C1(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__o211ai_1 _09042_ (.A1(_01658_),
    .A2(_01657_),
    .B1(_01562_),
    .C1(_01560_),
    .Y(_01660_));
 sky130_fd_sc_hd__o211ai_2 _09043_ (.A1(_01646_),
    .A2(_01585_),
    .B1(_01659_),
    .C1(_01660_),
    .Y(_01661_));
 sky130_fd_sc_hd__a211o_1 _09044_ (.A1(_01659_),
    .A2(_01660_),
    .B1(_01646_),
    .C1(_01585_),
    .X(_01662_));
 sky130_fd_sc_hd__a2bb2o_1 _09045_ (.A1_N(_01644_),
    .A2_N(_01645_),
    .B1(_01661_),
    .B2(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__or4bb_1 _09046_ (.A(_01644_),
    .B(_01645_),
    .C_N(_01661_),
    .D_N(_01662_),
    .X(_01664_));
 sky130_fd_sc_hd__o211a_2 _09047_ (.A1(_01566_),
    .A2(_01590_),
    .B1(_01663_),
    .C1(_01664_),
    .X(_01665_));
 sky130_fd_sc_hd__a211oi_1 _09048_ (.A1(_01664_),
    .A2(_01663_),
    .B1(_01590_),
    .C1(_01566_),
    .Y(_01666_));
 sky130_fd_sc_hd__or2b_1 _09049_ (.A(_01578_),
    .B_N(_01582_),
    .X(_01667_));
 sky130_fd_sc_hd__o31a_1 _09050_ (.A1(_01208_),
    .A2(_01579_),
    .A3(_01581_),
    .B1(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__a21oi_1 _09051_ (.A1(_01586_),
    .A2(_01588_),
    .B1(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__and3_1 _09052_ (.A(_01586_),
    .B(_01588_),
    .C(_01668_),
    .X(_01670_));
 sky130_fd_sc_hd__nor2_1 _09053_ (.A(_01669_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor3b_2 _09054_ (.A(_01665_),
    .B(_01666_),
    .C_N(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__o21ba_1 _09055_ (.A1(_01665_),
    .A2(_01666_),
    .B1_N(_01671_),
    .X(_01673_));
 sky130_fd_sc_hd__or2_1 _09056_ (.A(_01672_),
    .B(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__xnor2_1 _09057_ (.A(_01626_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__xnor2_2 _09058_ (.A(_01437_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__and3_1 _09059_ (.A(_01625_),
    .B(_01622_),
    .C(_01624_),
    .X(_01677_));
 sky130_fd_sc_hd__a21oi_1 _09060_ (.A1(_01625_),
    .A2(_01622_),
    .B1(_01624_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _09061_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand3_1 _09062_ (.A(_01601_),
    .B(_01598_),
    .C(_01600_),
    .Y(_01680_));
 sky130_fd_sc_hd__and4_1 _09063_ (.A(_01332_),
    .B(_02334_),
    .C(_00032_),
    .D(_04767_),
    .X(_01681_));
 sky130_fd_sc_hd__a22o_1 _09064_ (.A1(_02334_),
    .A2(_00032_),
    .B1(_06611_),
    .B2(_01332_),
    .X(_01682_));
 sky130_fd_sc_hd__and2b_1 _09065_ (.A_N(_01681_),
    .B(_01682_),
    .X(_01683_));
 sky130_fd_sc_hd__nand2_1 _09066_ (.A(_06545_),
    .B(_04649_),
    .Y(_01684_));
 sky130_fd_sc_hd__xnor2_1 _09067_ (.A(_01683_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__or3_1 _09068_ (.A(_01596_),
    .B(_01594_),
    .C(_01595_),
    .X(_01686_));
 sky130_fd_sc_hd__o21ai_1 _09069_ (.A1(_01596_),
    .A2(_01595_),
    .B1(_01594_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_06488_),
    .B(_06611_),
    .Y(_01688_));
 sky130_fd_sc_hd__a22oi_2 _09071_ (.A1(_06491_),
    .A2(_06602_),
    .B1(_06604_),
    .B2(_06492_),
    .Y(_01689_));
 sky130_fd_sc_hd__and4_1 _09072_ (.A(_06494_),
    .B(_00150_),
    .C(net10),
    .D(net11),
    .X(_01690_));
 sky130_fd_sc_hd__o21bai_1 _09073_ (.A1(_01688_),
    .A2(_01689_),
    .B1_N(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__a21o_1 _09074_ (.A1(_01686_),
    .A2(_01687_),
    .B1(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nand3_1 _09075_ (.A(_01686_),
    .B(_01691_),
    .C(_01687_),
    .Y(_01693_));
 sky130_fd_sc_hd__a21bo_1 _09076_ (.A1(_01685_),
    .A2(_01692_),
    .B1_N(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__a21o_1 _09077_ (.A1(_01601_),
    .A2(_01598_),
    .B1(_01600_),
    .X(_01695_));
 sky130_fd_sc_hd__nand3_2 _09078_ (.A(_01680_),
    .B(_01694_),
    .C(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__a31o_1 _09079_ (.A1(_06545_),
    .A2(_00059_),
    .A3(_01682_),
    .B1(_01681_),
    .X(_01697_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_02528_),
    .B(_00085_),
    .Y(_01698_));
 sky130_fd_sc_hd__and2b_1 _09081_ (.A_N(_01344_),
    .B(_01343_),
    .X(_01699_));
 sky130_fd_sc_hd__xnor2_1 _09082_ (.A(_01698_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__xor2_1 _09083_ (.A(_01697_),
    .B(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__nand2_4 _09084_ (.A(_02528_),
    .B(_00093_),
    .Y(_01702_));
 sky130_fd_sc_hd__a22oi_2 _09085_ (.A1(_06516_),
    .A2(_00098_),
    .B1(_00047_),
    .B2(_06520_),
    .Y(_01703_));
 sky130_fd_sc_hd__and4_1 _09086_ (.A(_02420_),
    .B(_06513_),
    .C(_00084_),
    .D(_04574_),
    .X(_01704_));
 sky130_fd_sc_hd__o21ba_1 _09087_ (.A1(_01702_),
    .A2(_01703_),
    .B1_N(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__xnor2_1 _09088_ (.A(_01701_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__a21o_1 _09089_ (.A1(_01680_),
    .A2(_01695_),
    .B1(_01694_),
    .X(_01707_));
 sky130_fd_sc_hd__nand3_1 _09090_ (.A(_01696_),
    .B(_01706_),
    .C(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__a21oi_2 _09091_ (.A1(_01605_),
    .A2(_01606_),
    .B1(_01607_),
    .Y(_01709_));
 sky130_fd_sc_hd__and3_1 _09092_ (.A(_01605_),
    .B(_01606_),
    .C(_01607_),
    .X(_01710_));
 sky130_fd_sc_hd__a211oi_4 _09093_ (.A1(_01696_),
    .A2(_01708_),
    .B1(_01709_),
    .C1(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__o2bb2a_1 _09094_ (.A1_N(_06680_),
    .A2_N(_04305_),
    .B1(_01366_),
    .B2(_01367_),
    .X(_01712_));
 sky130_fd_sc_hd__nor2_1 _09095_ (.A(_01368_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__and4_1 _09096_ (.A(net68),
    .B(net38),
    .C(net123),
    .D(net34),
    .X(_01714_));
 sky130_fd_sc_hd__nand2_1 _09097_ (.A(net122),
    .B(_00266_),
    .Y(_01715_));
 sky130_fd_sc_hd__a22oi_2 _09098_ (.A1(_02647_),
    .A2(_00592_),
    .B1(_00089_),
    .B2(_02582_),
    .Y(_01716_));
 sky130_fd_sc_hd__or3_1 _09099_ (.A(_01714_),
    .B(_01715_),
    .C(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__or2b_1 _09100_ (.A(_01714_),
    .B_N(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__and2_1 _09101_ (.A(_01713_),
    .B(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__xor2_1 _09102_ (.A(_01713_),
    .B(_01718_),
    .X(_01720_));
 sky130_fd_sc_hd__o2bb2a_1 _09103_ (.A1_N(_06610_),
    .A2_N(_04122_),
    .B1(_01416_),
    .B2(_01417_),
    .X(_01721_));
 sky130_fd_sc_hd__nor2_2 _09104_ (.A(_01418_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__and2_1 _09105_ (.A(_01720_),
    .B(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(_01697_),
    .B(_01700_),
    .Y(_01724_));
 sky130_fd_sc_hd__or2b_1 _09107_ (.A(_01705_),
    .B_N(_01701_),
    .X(_01725_));
 sky130_fd_sc_hd__xnor2_1 _09108_ (.A(_01373_),
    .B(_01378_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21o_1 _09109_ (.A1(_01724_),
    .A2(_01725_),
    .B1(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__nand3_1 _09110_ (.A(_01724_),
    .B(_01725_),
    .C(_01726_),
    .Y(_01728_));
 sky130_fd_sc_hd__o211a_1 _09111_ (.A1(_01719_),
    .A2(_01723_),
    .B1(_01727_),
    .C1(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__a211oi_2 _09112_ (.A1(_01727_),
    .A2(_01728_),
    .B1(_01719_),
    .C1(_01723_),
    .Y(_01730_));
 sky130_fd_sc_hd__o211a_1 _09113_ (.A1(_01710_),
    .A2(_01709_),
    .B1(_01708_),
    .C1(_01696_),
    .X(_01731_));
 sky130_fd_sc_hd__nor4_4 _09114_ (.A(_01711_),
    .B(_01729_),
    .C(_01730_),
    .D(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__a2bb2o_1 _09115_ (.A1_N(_01611_),
    .A2_N(_01613_),
    .B1(_01614_),
    .B2(_01381_),
    .X(_01733_));
 sky130_fd_sc_hd__or4b_2 _09116_ (.A(_01612_),
    .B(_01611_),
    .C(_01613_),
    .D_N(_01614_),
    .X(_01734_));
 sky130_fd_sc_hd__o211ai_2 _09117_ (.A1(_01711_),
    .A2(_01732_),
    .B1(_01733_),
    .C1(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__o211a_1 _09118_ (.A1(_01711_),
    .A2(_01732_),
    .B1(_01733_),
    .C1(_01734_),
    .X(_01736_));
 sky130_fd_sc_hd__xnor2_1 _09119_ (.A(_01427_),
    .B(_01428_),
    .Y(_01737_));
 sky130_fd_sc_hd__a22o_1 _09120_ (.A1(_00011_),
    .A2(_04111_),
    .B1(_00272_),
    .B2(_06631_),
    .X(_01738_));
 sky130_fd_sc_hd__and4_1 _09121_ (.A(_06631_),
    .B(_06630_),
    .C(_04111_),
    .D(_04176_),
    .X(_01739_));
 sky130_fd_sc_hd__a31o_1 _09122_ (.A1(_02851_),
    .A2(_04057_),
    .A3(_01738_),
    .B1(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__o2bb2a_1 _09123_ (.A1_N(_00221_),
    .A2_N(_03873_),
    .B1(_01424_),
    .B2(_01425_),
    .X(_01741_));
 sky130_fd_sc_hd__nor2_2 _09124_ (.A(_01426_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__or2_1 _09125_ (.A(_01740_),
    .B(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__and4_1 _09126_ (.A(_02905_),
    .B(_02970_),
    .C(_03884_),
    .D(_03971_),
    .X(_01744_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(_01740_),
    .B(_01742_),
    .Y(_01745_));
 sky130_fd_sc_hd__a21bo_1 _09128_ (.A1(_01743_),
    .A2(_01744_),
    .B1_N(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__or2b_1 _09129_ (.A(_01737_),
    .B_N(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(_03067_),
    .B(_03917_),
    .Y(_01748_));
 sky130_fd_sc_hd__xor2_1 _09131_ (.A(_01737_),
    .B(_01746_),
    .X(_01749_));
 sky130_fd_sc_hd__or2_1 _09132_ (.A(_01748_),
    .B(_01749_),
    .X(_01750_));
 sky130_fd_sc_hd__inv_2 _09133_ (.A(_01727_),
    .Y(_01751_));
 sky130_fd_sc_hd__a22o_1 _09134_ (.A1(_01431_),
    .A2(_01432_),
    .B1(_01433_),
    .B2(_01408_),
    .X(_01752_));
 sky130_fd_sc_hd__o211a_1 _09135_ (.A1(_01751_),
    .A2(_01729_),
    .B1(_01752_),
    .C1(_01434_),
    .X(_01753_));
 sky130_fd_sc_hd__a211oi_1 _09136_ (.A1(_01434_),
    .A2(_01752_),
    .B1(_01729_),
    .C1(_01751_),
    .Y(_01754_));
 sky130_fd_sc_hd__a211oi_1 _09137_ (.A1(_01747_),
    .A2(_01750_),
    .B1(_01753_),
    .C1(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__o211a_1 _09138_ (.A1(_01753_),
    .A2(_01754_),
    .B1(_01747_),
    .C1(_01750_),
    .X(_01756_));
 sky130_fd_sc_hd__a211o_1 _09139_ (.A1(_01734_),
    .A2(_01733_),
    .B1(_01732_),
    .C1(_01711_),
    .X(_01757_));
 sky130_fd_sc_hd__or4b_2 _09140_ (.A(_01736_),
    .B(_01755_),
    .C(_01756_),
    .D_N(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__o211a_1 _09141_ (.A1(_01415_),
    .A2(_01435_),
    .B1(_01434_),
    .C1(_01431_),
    .X(_01759_));
 sky130_fd_sc_hd__o2bb2a_1 _09142_ (.A1_N(_01618_),
    .A2_N(_01619_),
    .B1(_01759_),
    .B2(_01436_),
    .X(_01760_));
 sky130_fd_sc_hd__and4b_1 _09143_ (.A_N(_01436_),
    .B(_01618_),
    .C(_01619_),
    .D(_01620_),
    .X(_01761_));
 sky130_fd_sc_hd__a211oi_1 _09144_ (.A1(_01735_),
    .A2(_01758_),
    .B1(_01760_),
    .C1(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _09145_ (.A(_01753_),
    .B(_01755_),
    .Y(_01763_));
 sky130_fd_sc_hd__o211a_1 _09146_ (.A1(_01761_),
    .A2(_01760_),
    .B1(_01758_),
    .C1(_01735_),
    .X(_01764_));
 sky130_fd_sc_hd__or3_1 _09147_ (.A(_01762_),
    .B(_01763_),
    .C(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__and2b_1 _09148_ (.A_N(_01762_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_2 _09149_ (.A(_01679_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__o21ai_1 _09150_ (.A1(_01762_),
    .A2(_01764_),
    .B1(_01763_),
    .Y(_01768_));
 sky130_fd_sc_hd__a22oi_2 _09151_ (.A1(_00162_),
    .A2(_04638_),
    .B1(_00033_),
    .B2(_00164_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand2_1 _09152_ (.A(_06475_),
    .B(_04585_),
    .Y(_01770_));
 sky130_fd_sc_hd__and4_1 _09153_ (.A(_02291_),
    .B(_06548_),
    .C(_00030_),
    .D(_04703_),
    .X(_01771_));
 sky130_fd_sc_hd__o21ba_1 _09154_ (.A1(_01769_),
    .A2(_01770_),
    .B1_N(_01771_),
    .X(_01772_));
 sky130_fd_sc_hd__nor2_1 _09155_ (.A(_01704_),
    .B(_01703_),
    .Y(_01773_));
 sky130_fd_sc_hd__xnor2_1 _09156_ (.A(_01702_),
    .B(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__or2b_1 _09157_ (.A(_01772_),
    .B_N(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__and4_1 _09158_ (.A(net107),
    .B(net66),
    .C(_00082_),
    .D(net36),
    .X(_01776_));
 sky130_fd_sc_hd__nand2_1 _09159_ (.A(net106),
    .B(_00089_),
    .Y(_01777_));
 sky130_fd_sc_hd__a22oi_1 _09160_ (.A1(_02474_),
    .A2(_00082_),
    .B1(_00084_),
    .B2(_06564_),
    .Y(_01778_));
 sky130_fd_sc_hd__or3_1 _09161_ (.A(_01776_),
    .B(_01777_),
    .C(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__and2b_1 _09162_ (.A_N(_01776_),
    .B(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__xnor2_1 _09163_ (.A(_01772_),
    .B(_01774_),
    .Y(_01781_));
 sky130_fd_sc_hd__or2b_1 _09164_ (.A(_01780_),
    .B_N(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__xnor2_1 _09165_ (.A(_01720_),
    .B(_01722_),
    .Y(_01783_));
 sky130_fd_sc_hd__a21oi_2 _09166_ (.A1(_01775_),
    .A2(_01782_),
    .B1(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o21ai_1 _09167_ (.A1(_01714_),
    .A2(_01716_),
    .B1(_01715_),
    .Y(_01785_));
 sky130_fd_sc_hd__a22o_1 _09168_ (.A1(_06579_),
    .A2(_00266_),
    .B1(_00592_),
    .B2(_02582_),
    .X(_01786_));
 sky130_fd_sc_hd__and4_1 _09169_ (.A(_02582_),
    .B(_02647_),
    .C(_00266_),
    .D(_00592_),
    .X(_01787_));
 sky130_fd_sc_hd__a31o_1 _09170_ (.A1(_02723_),
    .A2(_04186_),
    .A3(_01786_),
    .B1(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__nand3_1 _09171_ (.A(_01717_),
    .B(_01785_),
    .C(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__a21o_1 _09172_ (.A1(_01717_),
    .A2(_01785_),
    .B1(_01788_),
    .X(_01790_));
 sky130_fd_sc_hd__nand2_1 _09173_ (.A(_02851_),
    .B(_04046_),
    .Y(_01791_));
 sky130_fd_sc_hd__and2b_1 _09174_ (.A_N(_01739_),
    .B(_01738_),
    .X(_01792_));
 sky130_fd_sc_hd__xnor2_1 _09175_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand3_1 _09176_ (.A(_01789_),
    .B(_01790_),
    .C(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__and3_1 _09177_ (.A(_01775_),
    .B(_01782_),
    .C(_01783_),
    .X(_01795_));
 sky130_fd_sc_hd__a211oi_2 _09178_ (.A1(_01789_),
    .A2(_01794_),
    .B1(_01784_),
    .C1(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__xor2_1 _09179_ (.A(_01748_),
    .B(_01749_),
    .X(_01797_));
 sky130_fd_sc_hd__o21a_1 _09180_ (.A1(_01784_),
    .A2(_01796_),
    .B1(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__nor3_1 _09181_ (.A(_01784_),
    .B(_01796_),
    .C(_01797_),
    .Y(_01799_));
 sky130_fd_sc_hd__a22oi_1 _09182_ (.A1(_02970_),
    .A2(_03895_),
    .B1(_03982_),
    .B2(_02916_),
    .Y(_01800_));
 sky130_fd_sc_hd__or2_1 _09183_ (.A(_01744_),
    .B(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__and4_1 _09184_ (.A(_00877_),
    .B(_00011_),
    .C(_06446_),
    .D(_04111_),
    .X(_01802_));
 sky130_fd_sc_hd__a22oi_1 _09185_ (.A1(_02808_),
    .A2(_06443_),
    .B1(_00303_),
    .B2(_02765_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _09186_ (.A(_01802_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__a31o_1 _09187_ (.A1(_02862_),
    .A2(_03993_),
    .A3(_01804_),
    .B1(_01802_),
    .X(_01805_));
 sky130_fd_sc_hd__and2b_1 _09188_ (.A_N(_01801_),
    .B(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__inv_2 _09189_ (.A(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _09190_ (.A(_01743_),
    .B(_01745_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor4_1 _09191_ (.A(_01798_),
    .B(_01799_),
    .C(_01807_),
    .D(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__or2_1 _09192_ (.A(_01798_),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__a2bb2o_1 _09193_ (.A1_N(_01755_),
    .A2_N(_01756_),
    .B1(_01757_),
    .B2(_01735_),
    .X(_01811_));
 sky130_fd_sc_hd__nand3_1 _09194_ (.A(_01693_),
    .B(_01685_),
    .C(_01692_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _09195_ (.A(_01771_),
    .B(_01769_),
    .Y(_01813_));
 sky130_fd_sc_hd__xnor2_1 _09196_ (.A(_01813_),
    .B(_01770_),
    .Y(_01814_));
 sky130_fd_sc_hd__or3_1 _09197_ (.A(_01690_),
    .B(_01688_),
    .C(_01689_),
    .X(_01815_));
 sky130_fd_sc_hd__o21ai_1 _09198_ (.A1(_01690_),
    .A2(_01689_),
    .B1(_01688_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(_06460_),
    .B(_04703_),
    .Y(_01817_));
 sky130_fd_sc_hd__a22oi_2 _09200_ (.A1(_06463_),
    .A2(_04767_),
    .B1(_06602_),
    .B2(_02107_),
    .Y(_01818_));
 sky130_fd_sc_hd__and4_1 _09201_ (.A(_06469_),
    .B(_02194_),
    .C(_04767_),
    .D(net10),
    .X(_01819_));
 sky130_fd_sc_hd__o21bai_1 _09202_ (.A1(_01817_),
    .A2(_01818_),
    .B1_N(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21o_1 _09203_ (.A1(_01815_),
    .A2(_01816_),
    .B1(_01820_),
    .X(_01821_));
 sky130_fd_sc_hd__nand3_1 _09204_ (.A(_01815_),
    .B(_01820_),
    .C(_01816_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21bo_1 _09205_ (.A1(_01814_),
    .A2(_01821_),
    .B1_N(_01822_),
    .X(_01823_));
 sky130_fd_sc_hd__a21o_1 _09206_ (.A1(_01693_),
    .A2(_01692_),
    .B1(_01685_),
    .X(_01824_));
 sky130_fd_sc_hd__nand3_2 _09207_ (.A(_01812_),
    .B(_01823_),
    .C(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__xnor2_1 _09208_ (.A(_01781_),
    .B(_01780_),
    .Y(_01826_));
 sky130_fd_sc_hd__a21o_1 _09209_ (.A1(_01812_),
    .A2(_01824_),
    .B1(_01823_),
    .X(_01827_));
 sky130_fd_sc_hd__nand3_1 _09210_ (.A(_01825_),
    .B(_01826_),
    .C(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__a21oi_1 _09211_ (.A1(_01696_),
    .A2(_01707_),
    .B1(_01706_),
    .Y(_01829_));
 sky130_fd_sc_hd__and3_1 _09212_ (.A(_01696_),
    .B(_01706_),
    .C(_01707_),
    .X(_01830_));
 sky130_fd_sc_hd__a211oi_2 _09213_ (.A1(_01825_),
    .A2(_01828_),
    .B1(_01829_),
    .C1(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__inv_2 _09214_ (.A(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__o211a_1 _09215_ (.A1(_01784_),
    .A2(_01795_),
    .B1(_01789_),
    .C1(_01794_),
    .X(_01833_));
 sky130_fd_sc_hd__o211a_1 _09216_ (.A1(_01830_),
    .A2(_01829_),
    .B1(_01828_),
    .C1(_01825_),
    .X(_01834_));
 sky130_fd_sc_hd__or4_2 _09217_ (.A(_01831_),
    .B(_01796_),
    .C(_01833_),
    .D(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__o22a_1 _09218_ (.A1(_01729_),
    .A2(_01730_),
    .B1(_01731_),
    .B2(_01711_),
    .X(_01836_));
 sky130_fd_sc_hd__a211oi_2 _09219_ (.A1(_01832_),
    .A2(_01835_),
    .B1(_01836_),
    .C1(_01732_),
    .Y(_01837_));
 sky130_fd_sc_hd__o22a_1 _09220_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01807_),
    .B2(_01808_),
    .X(_01838_));
 sky130_fd_sc_hd__o211a_1 _09221_ (.A1(_01732_),
    .A2(_01836_),
    .B1(_01835_),
    .C1(_01832_),
    .X(_01839_));
 sky130_fd_sc_hd__nor4_2 _09222_ (.A(_01837_),
    .B(_01809_),
    .C(_01838_),
    .D(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__a211o_1 _09223_ (.A1(_01758_),
    .A2(_01811_),
    .B1(_01840_),
    .C1(_01837_),
    .X(_01841_));
 sky130_fd_sc_hd__o211ai_1 _09224_ (.A1(_01837_),
    .A2(_01840_),
    .B1(_01811_),
    .C1(_01758_),
    .Y(_01842_));
 sky130_fd_sc_hd__a21bo_1 _09225_ (.A1(_01810_),
    .A2(_01841_),
    .B1_N(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__and3_1 _09226_ (.A(_01765_),
    .B(_01768_),
    .C(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__or3_1 _09227_ (.A(_01677_),
    .B(_01678_),
    .C(_01766_),
    .X(_01845_));
 sky130_fd_sc_hd__a21boi_1 _09228_ (.A1(_01767_),
    .A2(_01844_),
    .B1_N(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__xor2_2 _09229_ (.A(_01676_),
    .B(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__nor3_2 _09230_ (.A(_01626_),
    .B(_01672_),
    .C(_01673_),
    .Y(_01848_));
 sky130_fd_sc_hd__a211oi_2 _09231_ (.A1(_01625_),
    .A2(_01674_),
    .B1(_01848_),
    .C1(_01437_),
    .Y(_01849_));
 sky130_fd_sc_hd__or2_1 _09232_ (.A(_01848_),
    .B(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__and4bb_1 _09233_ (.A_N(_01644_),
    .B_N(_01645_),
    .C(_01661_),
    .D(_01662_),
    .X(_01851_));
 sky130_fd_sc_hd__and4bb_1 _09234_ (.A_N(_01631_),
    .B_N(_01632_),
    .C(_01640_),
    .D(_01641_),
    .X(_01852_));
 sky130_fd_sc_hd__a2bb2o_1 _09235_ (.A1_N(_01298_),
    .A2_N(_01299_),
    .B1(_01242_),
    .B2(_01300_),
    .X(_01853_));
 sky130_fd_sc_hd__or4bb_1 _09236_ (.A(_01298_),
    .B(_01299_),
    .C_N(_01242_),
    .D_N(_01300_),
    .X(_01854_));
 sky130_fd_sc_hd__o211a_1 _09237_ (.A1(_01631_),
    .A2(_01852_),
    .B1(_01853_),
    .C1(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__a211oi_1 _09238_ (.A1(_01854_),
    .A2(_01853_),
    .B1(_01852_),
    .C1(_01631_),
    .Y(_01856_));
 sky130_fd_sc_hd__inv_2 _09239_ (.A(_01658_),
    .Y(_01857_));
 sky130_fd_sc_hd__o21a_1 _09240_ (.A1(_01262_),
    .A2(_01264_),
    .B1(_01266_),
    .X(_01858_));
 sky130_fd_sc_hd__nor3_1 _09241_ (.A(_01262_),
    .B(_01264_),
    .C(_01266_),
    .Y(_01859_));
 sky130_fd_sc_hd__a211oi_2 _09242_ (.A1(_01638_),
    .A2(_01640_),
    .B1(_01858_),
    .C1(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__o211a_1 _09243_ (.A1(_01859_),
    .A2(_01858_),
    .B1(_01640_),
    .C1(_01638_),
    .X(_01861_));
 sky130_fd_sc_hd__a211oi_2 _09244_ (.A1(_01650_),
    .A2(_01857_),
    .B1(_01860_),
    .C1(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__o211a_1 _09245_ (.A1(_01860_),
    .A2(_01861_),
    .B1(_01650_),
    .C1(_01857_),
    .X(_01863_));
 sky130_fd_sc_hd__o22ai_2 _09246_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01862_),
    .B2(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__or4_4 _09247_ (.A(_01855_),
    .B(_01856_),
    .C(_01862_),
    .D(_01863_),
    .X(_01865_));
 sky130_fd_sc_hd__o211a_1 _09248_ (.A1(_01644_),
    .A2(_01851_),
    .B1(_01864_),
    .C1(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__a211oi_2 _09249_ (.A1(_01865_),
    .A2(_01864_),
    .B1(_01851_),
    .C1(_01644_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(_01659_),
    .B(_01661_),
    .Y(_01868_));
 sky130_fd_sc_hd__clkinv_2 _09251_ (.A(_01655_),
    .Y(_01869_));
 sky130_fd_sc_hd__or2_1 _09252_ (.A(_01203_),
    .B(_01211_),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_01203_),
    .B(_01211_),
    .Y(_01871_));
 sky130_fd_sc_hd__a2bb2o_1 _09254_ (.A1_N(_01653_),
    .A2_N(_01869_),
    .B1(_01870_),
    .B2(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__xnor2_1 _09255_ (.A(_01868_),
    .B(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__o21ai_2 _09256_ (.A1(_01866_),
    .A2(_01867_),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__or3_2 _09257_ (.A(_01866_),
    .B(_01867_),
    .C(_01873_),
    .X(_01875_));
 sky130_fd_sc_hd__o211ai_4 _09258_ (.A1(_01665_),
    .A2(_01672_),
    .B1(_01874_),
    .C1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a211o_1 _09259_ (.A1(_01875_),
    .A2(_01874_),
    .B1(_01672_),
    .C1(_01665_),
    .X(_01877_));
 sky130_fd_sc_hd__nand3_2 _09260_ (.A(_01669_),
    .B(_01876_),
    .C(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__a21o_1 _09261_ (.A1(_01876_),
    .A2(_01877_),
    .B1(_01669_),
    .X(_01879_));
 sky130_fd_sc_hd__and2_1 _09262_ (.A(_01878_),
    .B(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__xor2_2 _09263_ (.A(_01850_),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__nand3_1 _09264_ (.A(_01842_),
    .B(_01810_),
    .C(_01841_),
    .Y(_01882_));
 sky130_fd_sc_hd__a21o_1 _09265_ (.A1(_01842_),
    .A2(_01841_),
    .B1(_01810_),
    .X(_01883_));
 sky130_fd_sc_hd__o21ai_1 _09266_ (.A1(_01776_),
    .A2(_01778_),
    .B1(_01777_),
    .Y(_01884_));
 sky130_fd_sc_hd__a22oi_2 _09267_ (.A1(_06548_),
    .A2(_00035_),
    .B1(_04638_),
    .B2(_02291_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(net108),
    .B(_00098_),
    .Y(_01886_));
 sky130_fd_sc_hd__and4_1 _09269_ (.A(_06479_),
    .B(_06480_),
    .C(net6),
    .D(net7),
    .X(_01887_));
 sky130_fd_sc_hd__o21bai_1 _09270_ (.A1(_01885_),
    .A2(_01886_),
    .B1_N(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__a21o_1 _09271_ (.A1(_01779_),
    .A2(_01884_),
    .B1(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(_06564_),
    .B(_00082_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_2 _09273_ (.A(_02474_),
    .B(_00089_),
    .Y(_01891_));
 sky130_fd_sc_hd__xor2_1 _09274_ (.A(_01890_),
    .B(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__nor2_1 _09275_ (.A(_01890_),
    .B(_01891_),
    .Y(_01893_));
 sky130_fd_sc_hd__a31o_1 _09276_ (.A1(_02550_),
    .A2(_04316_),
    .A3(_01892_),
    .B1(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__and3_1 _09277_ (.A(_01779_),
    .B(_01888_),
    .C(_01884_),
    .X(_01895_));
 sky130_fd_sc_hd__a21o_1 _09278_ (.A1(_01889_),
    .A2(_01894_),
    .B1(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__a21o_1 _09279_ (.A1(_01789_),
    .A2(_01790_),
    .B1(_01793_),
    .X(_01897_));
 sky130_fd_sc_hd__nand3_1 _09280_ (.A(_01794_),
    .B(_01896_),
    .C(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__and4_1 _09281_ (.A(_06578_),
    .B(_06579_),
    .C(_00271_),
    .D(_04229_),
    .X(_01899_));
 sky130_fd_sc_hd__a22oi_2 _09282_ (.A1(_06583_),
    .A2(_00287_),
    .B1(_00267_),
    .B2(_02593_),
    .Y(_01900_));
 sky130_fd_sc_hd__and4bb_1 _09283_ (.A_N(_01899_),
    .B_N(_01900_),
    .C(_02712_),
    .D(_04111_),
    .X(_01901_));
 sky130_fd_sc_hd__nor2_1 _09284_ (.A(_01899_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_1 _09285_ (.A(_06593_),
    .B(_00272_),
    .Y(_01903_));
 sky130_fd_sc_hd__and2b_1 _09286_ (.A_N(_01787_),
    .B(_01786_),
    .X(_01904_));
 sky130_fd_sc_hd__xnor2_1 _09287_ (.A(_01903_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__and2b_1 _09288_ (.A_N(_01902_),
    .B(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(_01905_),
    .B(_01902_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(_06610_),
    .B(_03971_),
    .Y(_01908_));
 sky130_fd_sc_hd__xnor2_1 _09291_ (.A(_01908_),
    .B(_01804_),
    .Y(_01909_));
 sky130_fd_sc_hd__and2_1 _09292_ (.A(_01907_),
    .B(_01909_),
    .X(_01910_));
 sky130_fd_sc_hd__a21o_1 _09293_ (.A1(_01794_),
    .A2(_01897_),
    .B1(_01896_),
    .X(_01911_));
 sky130_fd_sc_hd__o211ai_1 _09294_ (.A1(_01906_),
    .A2(_01910_),
    .B1(_01898_),
    .C1(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__nand2_1 _09295_ (.A(_01898_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _09296_ (.A(_01744_),
    .B(_01806_),
    .Y(_01914_));
 sky130_fd_sc_hd__xor2_1 _09297_ (.A(_01808_),
    .B(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__a22o_1 _09298_ (.A1(_00011_),
    .A2(_03960_),
    .B1(_06446_),
    .B2(_00012_),
    .X(_01916_));
 sky130_fd_sc_hd__and4_1 _09299_ (.A(_06631_),
    .B(_06630_),
    .C(_06436_),
    .D(_06446_),
    .X(_01917_));
 sky130_fd_sc_hd__a31o_1 _09300_ (.A1(_02862_),
    .A2(_03906_),
    .A3(_01916_),
    .B1(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__and3_1 _09301_ (.A(_02916_),
    .B(_03917_),
    .C(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__xnor2_1 _09302_ (.A(_01805_),
    .B(_01801_),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_1 _09303_ (.A(_01919_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__xnor2_1 _09304_ (.A(_01913_),
    .B(_01915_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _09305_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__a21oi_1 _09306_ (.A1(_01913_),
    .A2(_01915_),
    .B1(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__o22a_1 _09307_ (.A1(_01809_),
    .A2(_01838_),
    .B1(_01839_),
    .B2(_01837_),
    .X(_01925_));
 sky130_fd_sc_hd__nand3_1 _09308_ (.A(_01822_),
    .B(_01814_),
    .C(_01821_),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _09309_ (.A(_01885_),
    .B(_01887_),
    .Y(_01927_));
 sky130_fd_sc_hd__xnor2_1 _09310_ (.A(_01927_),
    .B(_01886_),
    .Y(_01928_));
 sky130_fd_sc_hd__or3_1 _09311_ (.A(_01819_),
    .B(_01817_),
    .C(_01818_),
    .X(_01929_));
 sky130_fd_sc_hd__o21ai_1 _09312_ (.A1(_01819_),
    .A2(_01818_),
    .B1(_01817_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand2_1 _09313_ (.A(net111),
    .B(_00030_),
    .Y(_01931_));
 sky130_fd_sc_hd__a22oi_2 _09314_ (.A1(_00150_),
    .A2(_00032_),
    .B1(_04767_),
    .B2(_06469_),
    .Y(_01932_));
 sky130_fd_sc_hd__and4_1 _09315_ (.A(_02096_),
    .B(net116),
    .C(net8),
    .D(_04767_),
    .X(_01933_));
 sky130_fd_sc_hd__o21bai_1 _09316_ (.A1(_01931_),
    .A2(_01932_),
    .B1_N(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__a21o_1 _09317_ (.A1(_01929_),
    .A2(_01930_),
    .B1(_01934_),
    .X(_01935_));
 sky130_fd_sc_hd__nand3_1 _09318_ (.A(_01929_),
    .B(_01934_),
    .C(_01930_),
    .Y(_01936_));
 sky130_fd_sc_hd__a21bo_1 _09319_ (.A1(_01928_),
    .A2(_01935_),
    .B1_N(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__a21o_1 _09320_ (.A1(_01822_),
    .A2(_01821_),
    .B1(_01814_),
    .X(_01938_));
 sky130_fd_sc_hd__nand3_2 _09321_ (.A(_01926_),
    .B(_01937_),
    .C(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__or2b_1 _09322_ (.A(_01895_),
    .B_N(_01889_),
    .X(_01940_));
 sky130_fd_sc_hd__xnor2_1 _09323_ (.A(_01940_),
    .B(_01894_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21o_1 _09324_ (.A1(_01926_),
    .A2(_01938_),
    .B1(_01937_),
    .X(_01942_));
 sky130_fd_sc_hd__nand3_1 _09325_ (.A(_01939_),
    .B(_01941_),
    .C(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21oi_2 _09326_ (.A1(_01825_),
    .A2(_01827_),
    .B1(_01826_),
    .Y(_01944_));
 sky130_fd_sc_hd__and3_1 _09327_ (.A(_01825_),
    .B(_01826_),
    .C(_01827_),
    .X(_01945_));
 sky130_fd_sc_hd__a211oi_4 _09328_ (.A1(_01939_),
    .A2(_01943_),
    .B1(_01944_),
    .C1(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__a211o_1 _09329_ (.A1(_01898_),
    .A2(_01911_),
    .B1(_01906_),
    .C1(_01910_),
    .X(_01947_));
 sky130_fd_sc_hd__nand2_1 _09330_ (.A(_01912_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__o211a_1 _09331_ (.A1(_01945_),
    .A2(_01944_),
    .B1(_01943_),
    .C1(_01939_),
    .X(_01949_));
 sky130_fd_sc_hd__nor3_1 _09332_ (.A(_01946_),
    .B(_01948_),
    .C(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__o22ai_2 _09333_ (.A1(_01796_),
    .A2(_01833_),
    .B1(_01834_),
    .B2(_01831_),
    .Y(_01951_));
 sky130_fd_sc_hd__o211ai_2 _09334_ (.A1(_01946_),
    .A2(_01950_),
    .B1(_01951_),
    .C1(_01835_),
    .Y(_01952_));
 sky130_fd_sc_hd__xor2_1 _09335_ (.A(_01921_),
    .B(_01922_),
    .X(_01953_));
 sky130_fd_sc_hd__a211o_1 _09336_ (.A1(_01835_),
    .A2(_01951_),
    .B1(_01950_),
    .C1(_01946_),
    .X(_01954_));
 sky130_fd_sc_hd__nand3_1 _09337_ (.A(_01952_),
    .B(_01953_),
    .C(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__o211a_1 _09338_ (.A1(_01840_),
    .A2(_01925_),
    .B1(_01955_),
    .C1(_01952_),
    .X(_01956_));
 sky130_fd_sc_hd__a211oi_1 _09339_ (.A1(_01952_),
    .A2(_01955_),
    .B1(_01925_),
    .C1(_01840_),
    .Y(_01957_));
 sky130_fd_sc_hd__o21bai_1 _09340_ (.A1(_01924_),
    .A2(_01956_),
    .B1_N(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__and3_1 _09341_ (.A(_01882_),
    .B(_01883_),
    .C(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__a21o_1 _09342_ (.A1(_01765_),
    .A2(_01768_),
    .B1(_01843_),
    .X(_01960_));
 sky130_fd_sc_hd__a21o_1 _09343_ (.A1(_01959_),
    .A2(_01960_),
    .B1(_01844_),
    .X(_01961_));
 sky130_fd_sc_hd__xnor2_2 _09344_ (.A(_01767_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__and2b_1 _09345_ (.A_N(_01844_),
    .B(_01960_),
    .X(_01963_));
 sky130_fd_sc_hd__a21o_1 _09346_ (.A1(_01882_),
    .A2(_01883_),
    .B1(_01958_),
    .X(_01964_));
 sky130_fd_sc_hd__nand3_1 _09347_ (.A(_01936_),
    .B(_01928_),
    .C(_01935_),
    .Y(_01965_));
 sky130_fd_sc_hd__a22oi_1 _09348_ (.A1(_06548_),
    .A2(_04509_),
    .B1(_00035_),
    .B2(_02291_),
    .Y(_01966_));
 sky130_fd_sc_hd__and4_1 _09349_ (.A(_06479_),
    .B(_06480_),
    .C(_00084_),
    .D(_04574_),
    .X(_01967_));
 sky130_fd_sc_hd__nor2_1 _09350_ (.A(_01966_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(_06544_),
    .B(_04445_),
    .Y(_01969_));
 sky130_fd_sc_hd__xnor2_1 _09352_ (.A(_01968_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__or3_1 _09353_ (.A(_01933_),
    .B(_01931_),
    .C(_01932_),
    .X(_01971_));
 sky130_fd_sc_hd__o21ai_1 _09354_ (.A1(_01933_),
    .A2(_01932_),
    .B1(_01931_),
    .Y(_01972_));
 sky130_fd_sc_hd__nand2_1 _09355_ (.A(net111),
    .B(_04574_),
    .Y(_01973_));
 sky130_fd_sc_hd__a22oi_2 _09356_ (.A1(_06495_),
    .A2(net7),
    .B1(_00032_),
    .B2(_06494_),
    .Y(_01974_));
 sky130_fd_sc_hd__and4_1 _09357_ (.A(_02096_),
    .B(_02194_),
    .C(net7),
    .D(net8),
    .X(_01975_));
 sky130_fd_sc_hd__o21bai_1 _09358_ (.A1(_01973_),
    .A2(_01974_),
    .B1_N(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__a21o_1 _09359_ (.A1(_01971_),
    .A2(_01972_),
    .B1(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__nand3_1 _09360_ (.A(_01971_),
    .B(_01976_),
    .C(_01972_),
    .Y(_01978_));
 sky130_fd_sc_hd__a21bo_1 _09361_ (.A1(_01970_),
    .A2(_01977_),
    .B1_N(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__a21o_1 _09362_ (.A1(_01936_),
    .A2(_01935_),
    .B1(_01928_),
    .X(_01980_));
 sky130_fd_sc_hd__nand3_2 _09363_ (.A(_01965_),
    .B(_01979_),
    .C(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__o21ba_1 _09364_ (.A1(_01966_),
    .A2(_01969_),
    .B1_N(_01967_),
    .X(_01982_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_06663_),
    .B(_04305_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_1 _09366_ (.A(_01983_),
    .B(_01892_),
    .Y(_01984_));
 sky130_fd_sc_hd__xnor2_1 _09367_ (.A(_01982_),
    .B(_01984_),
    .Y(_01985_));
 sky130_fd_sc_hd__and2_1 _09368_ (.A(net106),
    .B(_04229_),
    .X(_01986_));
 sky130_fd_sc_hd__a22o_1 _09369_ (.A1(_02474_),
    .A2(_00592_),
    .B1(_00089_),
    .B2(_06564_),
    .X(_01987_));
 sky130_fd_sc_hd__nand2_2 _09370_ (.A(_02420_),
    .B(_00592_),
    .Y(_01988_));
 sky130_fd_sc_hd__o2bb2a_1 _09371_ (.A1_N(_01986_),
    .A2_N(_01987_),
    .B1(_01891_),
    .B2(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__xnor2_1 _09372_ (.A(_01985_),
    .B(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__a21o_1 _09373_ (.A1(_01965_),
    .A2(_01980_),
    .B1(_01979_),
    .X(_01991_));
 sky130_fd_sc_hd__nand3_1 _09374_ (.A(_01981_),
    .B(_01990_),
    .C(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__a21oi_1 _09375_ (.A1(_01939_),
    .A2(_01942_),
    .B1(_01941_),
    .Y(_01993_));
 sky130_fd_sc_hd__and3_1 _09376_ (.A(_01939_),
    .B(_01941_),
    .C(_01942_),
    .X(_01994_));
 sky130_fd_sc_hd__a211oi_2 _09377_ (.A1(_01981_),
    .A2(_01992_),
    .B1(_01993_),
    .C1(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__a211o_1 _09378_ (.A1(_01981_),
    .A2(_01992_),
    .B1(_01993_),
    .C1(_01994_),
    .X(_01996_));
 sky130_fd_sc_hd__and4_1 _09379_ (.A(net68),
    .B(net38),
    .C(net126),
    .D(net125),
    .X(_01997_));
 sky130_fd_sc_hd__a22oi_1 _09380_ (.A1(_06579_),
    .A2(_04100_),
    .B1(_00271_),
    .B2(_06578_),
    .Y(_01998_));
 sky130_fd_sc_hd__and4bb_1 _09381_ (.A_N(_01997_),
    .B_N(_01998_),
    .C(net122),
    .D(_04035_),
    .X(_01999_));
 sky130_fd_sc_hd__nor2_1 _09382_ (.A(_01997_),
    .B(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__o2bb2a_1 _09383_ (.A1_N(_06593_),
    .A2_N(_04111_),
    .B1(_01899_),
    .B2(_01900_),
    .X(_02001_));
 sky130_fd_sc_hd__nor2_1 _09384_ (.A(_01901_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__and2b_1 _09385_ (.A_N(_02000_),
    .B(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__xnor2_1 _09386_ (.A(_02002_),
    .B(_02000_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2_1 _09387_ (.A(_02851_),
    .B(_03884_),
    .Y(_02005_));
 sky130_fd_sc_hd__and2b_1 _09388_ (.A_N(_01917_),
    .B(_01916_),
    .X(_02006_));
 sky130_fd_sc_hd__xnor2_1 _09389_ (.A(_02005_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__and2_1 _09390_ (.A(_02004_),
    .B(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__or2b_1 _09391_ (.A(_01982_),
    .B_N(_01984_),
    .X(_02009_));
 sky130_fd_sc_hd__or2b_1 _09392_ (.A(_01989_),
    .B_N(_01985_),
    .X(_02010_));
 sky130_fd_sc_hd__xnor2_1 _09393_ (.A(_01907_),
    .B(_01909_),
    .Y(_02011_));
 sky130_fd_sc_hd__a21o_1 _09394_ (.A1(_02009_),
    .A2(_02010_),
    .B1(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__nand3_1 _09395_ (.A(_02009_),
    .B(_02010_),
    .C(_02011_),
    .Y(_02013_));
 sky130_fd_sc_hd__o211ai_2 _09396_ (.A1(_02003_),
    .A2(_02008_),
    .B1(_02012_),
    .C1(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__a211o_1 _09397_ (.A1(_02012_),
    .A2(_02013_),
    .B1(_02003_),
    .C1(_02008_),
    .X(_02015_));
 sky130_fd_sc_hd__o211ai_1 _09398_ (.A1(_01994_),
    .A2(_01993_),
    .B1(_01992_),
    .C1(_01981_),
    .Y(_02016_));
 sky130_fd_sc_hd__and4_1 _09399_ (.A(_01996_),
    .B(_02014_),
    .C(_02015_),
    .D(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__o21ai_2 _09400_ (.A1(_01946_),
    .A2(_01949_),
    .B1(_01948_),
    .Y(_02018_));
 sky130_fd_sc_hd__or3_1 _09401_ (.A(_01946_),
    .B(_01948_),
    .C(_01949_),
    .X(_02019_));
 sky130_fd_sc_hd__o211ai_4 _09402_ (.A1(_01995_),
    .A2(_02017_),
    .B1(_02018_),
    .C1(_02019_),
    .Y(_02021_));
 sky130_fd_sc_hd__or2_1 _09403_ (.A(_01919_),
    .B(_01920_),
    .X(_02022_));
 sky130_fd_sc_hd__nand2_1 _09404_ (.A(_01921_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__a21oi_1 _09405_ (.A1(_02012_),
    .A2(_02014_),
    .B1(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__and3_1 _09406_ (.A(_02012_),
    .B(_02014_),
    .C(_02023_),
    .X(_02025_));
 sky130_fd_sc_hd__nor2_1 _09407_ (.A(_02024_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__a211o_1 _09408_ (.A1(_02019_),
    .A2(_02018_),
    .B1(_02017_),
    .C1(_01995_),
    .X(_02027_));
 sky130_fd_sc_hd__nand3_2 _09409_ (.A(_02021_),
    .B(_02026_),
    .C(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__a21oi_1 _09410_ (.A1(_01952_),
    .A2(_01954_),
    .B1(_01953_),
    .Y(_02029_));
 sky130_fd_sc_hd__and3_1 _09411_ (.A(_01952_),
    .B(_01953_),
    .C(_01954_),
    .X(_02030_));
 sky130_fd_sc_hd__a211oi_2 _09412_ (.A1(_02021_),
    .A2(_02028_),
    .B1(_02029_),
    .C1(_02030_),
    .Y(_02032_));
 sky130_fd_sc_hd__o211a_1 _09413_ (.A1(_02030_),
    .A2(_02029_),
    .B1(_02028_),
    .C1(_02021_),
    .X(_02033_));
 sky130_fd_sc_hd__nor3b_2 _09414_ (.A(_02032_),
    .B(_02033_),
    .C_N(_02024_),
    .Y(_02034_));
 sky130_fd_sc_hd__or3_1 _09415_ (.A(_01957_),
    .B(_01924_),
    .C(_01956_),
    .X(_02035_));
 sky130_fd_sc_hd__o21ai_1 _09416_ (.A1(_01957_),
    .A2(_01956_),
    .B1(_01924_),
    .Y(_02036_));
 sky130_fd_sc_hd__o211a_1 _09417_ (.A1(_02032_),
    .A2(_02034_),
    .B1(_02035_),
    .C1(_02036_),
    .X(_02037_));
 sky130_fd_sc_hd__a21oi_1 _09418_ (.A1(_01964_),
    .A2(_02037_),
    .B1(_01959_),
    .Y(_02038_));
 sky130_fd_sc_hd__xnor2_1 _09419_ (.A(_01963_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__and2b_1 _09420_ (.A_N(_01962_),
    .B(_02039_),
    .X(_02040_));
 sky130_fd_sc_hd__and3_1 _09421_ (.A(_01847_),
    .B(_01881_),
    .C(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__and4_1 _09422_ (.A(_06479_),
    .B(_06480_),
    .C(net34),
    .D(_00082_),
    .X(_02043_));
 sky130_fd_sc_hd__a22oi_1 _09423_ (.A1(_06504_),
    .A2(_00072_),
    .B1(_04434_),
    .B2(_06503_),
    .Y(_02044_));
 sky130_fd_sc_hd__and4bb_1 _09424_ (.A_N(_02043_),
    .B_N(_02044_),
    .C(_06544_),
    .D(_00074_),
    .X(_02045_));
 sky130_fd_sc_hd__nor2_1 _09425_ (.A(_02043_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__nand2_1 _09426_ (.A(_06663_),
    .B(_04176_),
    .Y(_02047_));
 sky130_fd_sc_hd__and4_1 _09427_ (.A(_06519_),
    .B(_06515_),
    .C(net124),
    .D(net123),
    .X(_02048_));
 sky130_fd_sc_hd__a22o_1 _09428_ (.A1(_06515_),
    .A2(net124),
    .B1(net123),
    .B2(_06519_),
    .X(_02049_));
 sky130_fd_sc_hd__and2b_1 _09429_ (.A_N(_02048_),
    .B(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__xnor2_1 _09430_ (.A(_02047_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__or2b_1 _09431_ (.A(_02046_),
    .B_N(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__and4_1 _09432_ (.A(_02442_),
    .B(_02496_),
    .C(_00272_),
    .D(_00301_),
    .X(_02054_));
 sky130_fd_sc_hd__nand4_1 _09433_ (.A(_06520_),
    .B(_06513_),
    .C(_00271_),
    .D(_04229_),
    .Y(_02055_));
 sky130_fd_sc_hd__a22o_1 _09434_ (.A1(_02474_),
    .A2(_04165_),
    .B1(_00266_),
    .B2(_06564_),
    .X(_02056_));
 sky130_fd_sc_hd__and4_1 _09435_ (.A(_06663_),
    .B(_06433_),
    .C(_02055_),
    .D(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__nor2_1 _09436_ (.A(_02054_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_1 _09437_ (.A(_02046_),
    .B(_02051_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2b_1 _09438_ (.A(_02058_),
    .B_N(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__o2bb2a_1 _09439_ (.A1_N(_06680_),
    .A2_N(_04035_),
    .B1(_01997_),
    .B2(_01998_),
    .X(_02061_));
 sky130_fd_sc_hd__nor2_1 _09440_ (.A(_01999_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__and4_1 _09441_ (.A(net68),
    .B(net38),
    .C(net127),
    .D(net126),
    .X(_02063_));
 sky130_fd_sc_hd__a22oi_2 _09442_ (.A1(_06579_),
    .A2(net127),
    .B1(_06431_),
    .B2(_06578_),
    .Y(_02065_));
 sky130_fd_sc_hd__and4bb_1 _09443_ (.A_N(_02063_),
    .B_N(_02065_),
    .C(net122),
    .D(_06436_),
    .X(_02066_));
 sky130_fd_sc_hd__nor2_1 _09444_ (.A(_02063_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__xnor2_1 _09445_ (.A(_02062_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__and4_2 _09446_ (.A(_02754_),
    .B(_02797_),
    .C(net115),
    .D(net132),
    .X(_02069_));
 sky130_fd_sc_hd__a22oi_1 _09447_ (.A1(_06630_),
    .A2(net115),
    .B1(_03960_),
    .B2(_06631_),
    .Y(_02070_));
 sky130_fd_sc_hd__or2_1 _09448_ (.A(_02069_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__inv_2 _09449_ (.A(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__xnor2_1 _09450_ (.A(_02068_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__a21oi_2 _09451_ (.A1(_02052_),
    .A2(_02060_),
    .B1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__o2bb2a_1 _09452_ (.A1_N(_06620_),
    .A2_N(_06437_),
    .B1(_02063_),
    .B2(_02065_),
    .X(_02076_));
 sky130_fd_sc_hd__and4_1 _09453_ (.A(_02593_),
    .B(_06583_),
    .C(_06436_),
    .D(_06430_),
    .X(_02077_));
 sky130_fd_sc_hd__a22oi_4 _09454_ (.A1(_06682_),
    .A2(_06436_),
    .B1(_06446_),
    .B2(_00000_),
    .Y(_02078_));
 sky130_fd_sc_hd__and4bb_1 _09455_ (.A_N(_02077_),
    .B_N(_02078_),
    .C(_06620_),
    .D(_03873_),
    .X(_02079_));
 sky130_fd_sc_hd__nor2_1 _09456_ (.A(_02077_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__or3_1 _09457_ (.A(_02066_),
    .B(_02076_),
    .C(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__nand2_1 _09458_ (.A(_02765_),
    .B(_03895_),
    .Y(_02082_));
 sky130_fd_sc_hd__nor2_1 _09459_ (.A(_02066_),
    .B(_02076_),
    .Y(_02083_));
 sky130_fd_sc_hd__xnor2_1 _09460_ (.A(_02083_),
    .B(_02080_),
    .Y(_02084_));
 sky130_fd_sc_hd__or2b_1 _09461_ (.A(_02082_),
    .B_N(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__and3_1 _09462_ (.A(_02052_),
    .B(_02060_),
    .C(_02073_),
    .X(_02086_));
 sky130_fd_sc_hd__a211oi_2 _09463_ (.A1(_02081_),
    .A2(_02085_),
    .B1(_02074_),
    .C1(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__o21ai_2 _09464_ (.A1(_02074_),
    .A2(_02087_),
    .B1(_02069_),
    .Y(_02088_));
 sky130_fd_sc_hd__or3_1 _09465_ (.A(_02069_),
    .B(_02074_),
    .C(_02087_),
    .X(_02089_));
 sky130_fd_sc_hd__and2_1 _09466_ (.A(_02088_),
    .B(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_02248_),
    .B(_00098_),
    .Y(_02091_));
 sky130_fd_sc_hd__and4_1 _09468_ (.A(_06494_),
    .B(_00150_),
    .C(net6),
    .D(net7),
    .X(_02092_));
 sky130_fd_sc_hd__a22oi_2 _09469_ (.A1(_02205_),
    .A2(_00035_),
    .B1(_00030_),
    .B2(_06534_),
    .Y(_02093_));
 sky130_fd_sc_hd__or3_1 _09470_ (.A(_02091_),
    .B(_02092_),
    .C(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__o21ai_1 _09471_ (.A1(_02092_),
    .A2(_02093_),
    .B1(_02091_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _09472_ (.A(_06488_),
    .B(_04434_),
    .Y(_02097_));
 sky130_fd_sc_hd__a22oi_2 _09473_ (.A1(_06491_),
    .A2(_04509_),
    .B1(_00035_),
    .B2(_06534_),
    .Y(_02098_));
 sky130_fd_sc_hd__and4_1 _09474_ (.A(_06494_),
    .B(_06495_),
    .C(_00084_),
    .D(_04574_),
    .X(_02099_));
 sky130_fd_sc_hd__o21bai_1 _09475_ (.A1(_02097_),
    .A2(_02098_),
    .B1_N(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__a21o_1 _09476_ (.A1(_02094_),
    .A2(_02095_),
    .B1(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__o2bb2a_1 _09477_ (.A1_N(_06545_),
    .A2_N(_00259_),
    .B1(_02043_),
    .B2(_02044_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_02045_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand3_1 _09479_ (.A(_02100_),
    .B(_02094_),
    .C(_02095_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21bo_1 _09480_ (.A1(_02101_),
    .A2(_02103_),
    .B1_N(_02104_),
    .X(_02105_));
 sky130_fd_sc_hd__or3_1 _09481_ (.A(_01975_),
    .B(_01973_),
    .C(_01974_),
    .X(_02106_));
 sky130_fd_sc_hd__o21bai_1 _09482_ (.A1(_02091_),
    .A2(_02093_),
    .B1_N(_02092_),
    .Y(_02108_));
 sky130_fd_sc_hd__o21ai_1 _09483_ (.A1(_01975_),
    .A2(_01974_),
    .B1(_01973_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand3_1 _09484_ (.A(_02106_),
    .B(_02108_),
    .C(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__a21o_1 _09485_ (.A1(_02106_),
    .A2(_02109_),
    .B1(_02108_),
    .X(_02111_));
 sky130_fd_sc_hd__nand2_1 _09486_ (.A(_06544_),
    .B(_04358_),
    .Y(_02112_));
 sky130_fd_sc_hd__a22oi_1 _09487_ (.A1(_06548_),
    .A2(_04434_),
    .B1(_00098_),
    .B2(_02291_),
    .Y(_02113_));
 sky130_fd_sc_hd__and4_1 _09488_ (.A(_01332_),
    .B(_02334_),
    .C(_00082_),
    .D(_00084_),
    .X(_02114_));
 sky130_fd_sc_hd__nor2_1 _09489_ (.A(_02113_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__xnor2_1 _09490_ (.A(_02112_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand3_1 _09491_ (.A(_02110_),
    .B(_02111_),
    .C(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21o_1 _09492_ (.A1(_02110_),
    .A2(_02111_),
    .B1(_02116_),
    .X(_02119_));
 sky130_fd_sc_hd__nand3_2 _09493_ (.A(_02105_),
    .B(_02117_),
    .C(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21o_1 _09494_ (.A1(_02117_),
    .A2(_02119_),
    .B1(_02105_),
    .X(_02121_));
 sky130_fd_sc_hd__xnor2_1 _09495_ (.A(_02058_),
    .B(_02059_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand3_1 _09496_ (.A(_02120_),
    .B(_02121_),
    .C(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_01978_),
    .B(_01970_),
    .C(_01977_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21bo_1 _09498_ (.A1(_02111_),
    .A2(_02116_),
    .B1_N(_02110_),
    .X(_02125_));
 sky130_fd_sc_hd__a21o_1 _09499_ (.A1(_01978_),
    .A2(_01977_),
    .B1(_01970_),
    .X(_02126_));
 sky130_fd_sc_hd__nand3_2 _09500_ (.A(_02124_),
    .B(_02125_),
    .C(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__a21o_1 _09501_ (.A1(_02124_),
    .A2(_02126_),
    .B1(_02125_),
    .X(_02128_));
 sky130_fd_sc_hd__a31o_1 _09502_ (.A1(_02539_),
    .A2(_04186_),
    .A3(_02049_),
    .B1(_02048_),
    .X(_02130_));
 sky130_fd_sc_hd__o21ba_1 _09503_ (.A1(_02112_),
    .A2(_02113_),
    .B1_N(_02114_),
    .X(_02131_));
 sky130_fd_sc_hd__o21ai_1 _09504_ (.A1(_01891_),
    .A2(_01988_),
    .B1(_01987_),
    .Y(_02132_));
 sky130_fd_sc_hd__xnor2_1 _09505_ (.A(_01986_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__xnor2_1 _09506_ (.A(_02131_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__xor2_1 _09507_ (.A(_02130_),
    .B(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__and3_1 _09508_ (.A(_02127_),
    .B(_02128_),
    .C(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__a21oi_1 _09509_ (.A1(_02127_),
    .A2(_02128_),
    .B1(_02135_),
    .Y(_02137_));
 sky130_fd_sc_hd__a211o_1 _09510_ (.A1(_02120_),
    .A2(_02123_),
    .B1(_02136_),
    .C1(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__a211oi_1 _09511_ (.A1(_02120_),
    .A2(_02123_),
    .B1(_02136_),
    .C1(_02137_),
    .Y(_02139_));
 sky130_fd_sc_hd__o211a_1 _09512_ (.A1(_02136_),
    .A2(_02137_),
    .B1(_02120_),
    .C1(_02123_),
    .X(_02141_));
 sky130_fd_sc_hd__o211a_1 _09513_ (.A1(_02074_),
    .A2(_02086_),
    .B1(_02081_),
    .C1(_02085_),
    .X(_02142_));
 sky130_fd_sc_hd__or4_2 _09514_ (.A(_02087_),
    .B(_02139_),
    .C(_02141_),
    .D(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__nand3_1 _09515_ (.A(_02127_),
    .B(_02128_),
    .C(_02135_),
    .Y(_02144_));
 sky130_fd_sc_hd__a21oi_1 _09516_ (.A1(_01981_),
    .A2(_01991_),
    .B1(_01990_),
    .Y(_02145_));
 sky130_fd_sc_hd__and3_1 _09517_ (.A(_01981_),
    .B(_01990_),
    .C(_01991_),
    .X(_02146_));
 sky130_fd_sc_hd__a211oi_2 _09518_ (.A1(_02127_),
    .A2(_02144_),
    .B1(_02145_),
    .C1(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__o211a_1 _09519_ (.A1(_02146_),
    .A2(_02145_),
    .B1(_02144_),
    .C1(_02127_),
    .X(_02148_));
 sky130_fd_sc_hd__or2b_1 _09520_ (.A(_02131_),
    .B_N(_02133_),
    .X(_02149_));
 sky130_fd_sc_hd__nand2_1 _09521_ (.A(_02130_),
    .B(_02134_),
    .Y(_02150_));
 sky130_fd_sc_hd__xnor2_1 _09522_ (.A(_02004_),
    .B(_02007_),
    .Y(_02152_));
 sky130_fd_sc_hd__a21o_1 _09523_ (.A1(_02149_),
    .A2(_02150_),
    .B1(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__nand3_1 _09524_ (.A(_02149_),
    .B(_02150_),
    .C(_02152_),
    .Y(_02154_));
 sky130_fd_sc_hd__or3_1 _09525_ (.A(_01999_),
    .B(_02061_),
    .C(_02067_),
    .X(_02155_));
 sky130_fd_sc_hd__a21bo_1 _09526_ (.A1(_02068_),
    .A2(_02072_),
    .B1_N(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__nand3_1 _09527_ (.A(_02153_),
    .B(_02154_),
    .C(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__a21o_1 _09528_ (.A1(_02153_),
    .A2(_02154_),
    .B1(_02156_),
    .X(_02158_));
 sky130_fd_sc_hd__and4bb_1 _09529_ (.A_N(_02147_),
    .B_N(_02148_),
    .C(_02157_),
    .D(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__a2bb2oi_1 _09530_ (.A1_N(_02147_),
    .A2_N(_02148_),
    .B1(_02157_),
    .B2(_02158_),
    .Y(_02160_));
 sky130_fd_sc_hd__a211o_1 _09531_ (.A1(_02138_),
    .A2(_02143_),
    .B1(_02159_),
    .C1(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__o211ai_1 _09532_ (.A1(_02159_),
    .A2(_02160_),
    .B1(_02138_),
    .C1(_02143_),
    .Y(_02163_));
 sky130_fd_sc_hd__and3_1 _09533_ (.A(_02090_),
    .B(_02161_),
    .C(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__a21oi_1 _09534_ (.A1(_02161_),
    .A2(_02163_),
    .B1(_02090_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _09535_ (.A(_02164_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__o2bb2a_1 _09536_ (.A1_N(_06620_),
    .A2_N(_03873_),
    .B1(_02077_),
    .B2(_02078_),
    .X(_02167_));
 sky130_fd_sc_hd__nor2_1 _09537_ (.A(_02079_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__and4_1 _09538_ (.A(_02604_),
    .B(_02669_),
    .C(_03873_),
    .D(_03971_),
    .X(_02169_));
 sky130_fd_sc_hd__and2_1 _09539_ (.A(_02168_),
    .B(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _09540_ (.A1(_06504_),
    .A2(_04294_),
    .B1(_00072_),
    .B2(_06503_),
    .X(_02171_));
 sky130_fd_sc_hd__and4_1 _09541_ (.A(_01332_),
    .B(_02334_),
    .C(_00592_),
    .D(_00089_),
    .X(_02172_));
 sky130_fd_sc_hd__a31o_1 _09542_ (.A1(_06545_),
    .A2(_04251_),
    .A3(_02171_),
    .B1(_02172_),
    .X(_02174_));
 sky130_fd_sc_hd__a22o_1 _09543_ (.A1(_02528_),
    .A2(_04111_),
    .B1(_02055_),
    .B2(_02056_),
    .X(_02175_));
 sky130_fd_sc_hd__and2b_1 _09544_ (.A_N(_02057_),
    .B(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__xor2_1 _09545_ (.A(_02174_),
    .B(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__a22o_1 _09546_ (.A1(_06513_),
    .A2(_04100_),
    .B1(_04165_),
    .B2(_02420_),
    .X(_02178_));
 sky130_fd_sc_hd__and4_1 _09547_ (.A(_06564_),
    .B(_02474_),
    .C(_04100_),
    .D(_04165_),
    .X(_02179_));
 sky130_fd_sc_hd__a31oi_4 _09548_ (.A1(_02550_),
    .A2(_04057_),
    .A3(_02178_),
    .B1(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__inv_2 _09549_ (.A(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__and2_1 _09550_ (.A(_02174_),
    .B(_02176_),
    .X(_02182_));
 sky130_fd_sc_hd__a21oi_1 _09551_ (.A1(_02177_),
    .A2(_02181_),
    .B1(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__xnor2_1 _09552_ (.A(_02082_),
    .B(_02084_),
    .Y(_02184_));
 sky130_fd_sc_hd__xnor2_1 _09553_ (.A(_02183_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__and2b_1 _09554_ (.A_N(_02183_),
    .B(_02184_),
    .X(_02186_));
 sky130_fd_sc_hd__a21o_1 _09555_ (.A1(_02170_),
    .A2(_02185_),
    .B1(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__o22ai_1 _09556_ (.A1(_02139_),
    .A2(_02141_),
    .B1(_02142_),
    .B2(_02087_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand3_1 _09557_ (.A(_02104_),
    .B(_02101_),
    .C(_02103_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21o_1 _09558_ (.A1(_02104_),
    .A2(_02101_),
    .B1(_02103_),
    .X(_02190_));
 sky130_fd_sc_hd__and2b_1 _09559_ (.A_N(_02172_),
    .B(_02171_),
    .X(_02191_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_02377_),
    .B(_00301_),
    .Y(_02192_));
 sky130_fd_sc_hd__xnor2_1 _09561_ (.A(_02191_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__or3_1 _09562_ (.A(_02099_),
    .B(_02097_),
    .C(_02098_),
    .X(_02195_));
 sky130_fd_sc_hd__o21ai_1 _09563_ (.A1(_02099_),
    .A2(_02098_),
    .B1(_02097_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _09564_ (.A(_06488_),
    .B(_00072_),
    .Y(_02197_));
 sky130_fd_sc_hd__a22oi_2 _09565_ (.A1(_06491_),
    .A2(_04434_),
    .B1(_04509_),
    .B2(_06492_),
    .Y(_02198_));
 sky130_fd_sc_hd__and4_1 _09566_ (.A(_06494_),
    .B(_06495_),
    .C(_00082_),
    .D(_00084_),
    .X(_02199_));
 sky130_fd_sc_hd__o21bai_1 _09567_ (.A1(_02197_),
    .A2(_02198_),
    .B1_N(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__a21o_1 _09568_ (.A1(_02195_),
    .A2(_02196_),
    .B1(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__nand3_1 _09569_ (.A(_02195_),
    .B(_02196_),
    .C(_02200_),
    .Y(_02202_));
 sky130_fd_sc_hd__a21bo_1 _09570_ (.A1(_02193_),
    .A2(_02201_),
    .B1_N(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__nand3_2 _09571_ (.A(_02189_),
    .B(_02190_),
    .C(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__xnor2_1 _09572_ (.A(_02177_),
    .B(_02180_),
    .Y(_02206_));
 sky130_fd_sc_hd__a21o_1 _09573_ (.A1(_02189_),
    .A2(_02190_),
    .B1(_02203_),
    .X(_02207_));
 sky130_fd_sc_hd__nand3_2 _09574_ (.A(_02204_),
    .B(_02206_),
    .C(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__and3_1 _09575_ (.A(_02120_),
    .B(_02121_),
    .C(_02122_),
    .X(_02209_));
 sky130_fd_sc_hd__a21oi_1 _09576_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_02122_),
    .Y(_02210_));
 sky130_fd_sc_hd__a211oi_2 _09577_ (.A1(_02204_),
    .A2(_02208_),
    .B1(_02209_),
    .C1(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__xnor2_1 _09578_ (.A(_02170_),
    .B(_02185_),
    .Y(_02212_));
 sky130_fd_sc_hd__o211a_1 _09579_ (.A1(_02209_),
    .A2(_02210_),
    .B1(_02204_),
    .C1(_02208_),
    .X(_02213_));
 sky130_fd_sc_hd__nor3_1 _09580_ (.A(_02211_),
    .B(_02212_),
    .C(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__a211o_1 _09581_ (.A1(_02143_),
    .A2(_02188_),
    .B1(_02211_),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__o211a_1 _09582_ (.A1(_02211_),
    .A2(_02214_),
    .B1(_02143_),
    .C1(_02188_),
    .X(_02217_));
 sky130_fd_sc_hd__a21o_1 _09583_ (.A1(_02187_),
    .A2(_02215_),
    .B1(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__xnor2_1 _09584_ (.A(_02166_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__a22o_1 _09585_ (.A1(_02334_),
    .A2(_00266_),
    .B1(_04294_),
    .B2(_01332_),
    .X(_02220_));
 sky130_fd_sc_hd__and4_1 _09586_ (.A(_01332_),
    .B(_06480_),
    .C(_00266_),
    .D(_00592_),
    .X(_02221_));
 sky130_fd_sc_hd__a31o_1 _09587_ (.A1(_06545_),
    .A2(_04186_),
    .A3(_02220_),
    .B1(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__nand2_1 _09588_ (.A(_06560_),
    .B(_06443_),
    .Y(_02223_));
 sky130_fd_sc_hd__and2b_1 _09589_ (.A_N(_02179_),
    .B(_02178_),
    .X(_02224_));
 sky130_fd_sc_hd__xnor2_1 _09590_ (.A(_02223_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(_02222_),
    .B(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _09592_ (.A(_06560_),
    .B(_03960_),
    .Y(_02228_));
 sky130_fd_sc_hd__buf_4 _09593_ (.A(_06513_),
    .X(_02229_));
 sky130_fd_sc_hd__a22oi_2 _09594_ (.A1(_02229_),
    .A2(_04035_),
    .B1(_06433_),
    .B2(_02431_),
    .Y(_02230_));
 sky130_fd_sc_hd__and4_1 _09595_ (.A(_06520_),
    .B(_06516_),
    .C(_06430_),
    .D(_06431_),
    .X(_02231_));
 sky130_fd_sc_hd__o21ba_1 _09596_ (.A1(_02228_),
    .A2(_02230_),
    .B1_N(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__xor2_1 _09597_ (.A(_02222_),
    .B(_02225_),
    .X(_02233_));
 sky130_fd_sc_hd__or2b_1 _09598_ (.A(_02232_),
    .B_N(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__nor2_1 _09599_ (.A(_02168_),
    .B(_02169_),
    .Y(_02235_));
 sky130_fd_sc_hd__or2_1 _09600_ (.A(_02170_),
    .B(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__a21oi_1 _09601_ (.A1(_02226_),
    .A2(_02234_),
    .B1(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand3_1 _09602_ (.A(_02202_),
    .B(_02193_),
    .C(_02201_),
    .Y(_02238_));
 sky130_fd_sc_hd__a21o_1 _09603_ (.A1(_02202_),
    .A2(_02201_),
    .B1(_02193_),
    .X(_02239_));
 sky130_fd_sc_hd__and2b_1 _09604_ (.A_N(_02221_),
    .B(_02220_),
    .X(_02240_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_02377_),
    .B(_00272_),
    .Y(_02241_));
 sky130_fd_sc_hd__xnor2_1 _09606_ (.A(_02240_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__or3_1 _09607_ (.A(_02199_),
    .B(_02197_),
    .C(_02198_),
    .X(_02243_));
 sky130_fd_sc_hd__o21ai_1 _09608_ (.A1(_02199_),
    .A2(_02198_),
    .B1(_02197_),
    .Y(_02244_));
 sky130_fd_sc_hd__and2_1 _09609_ (.A(_06488_),
    .B(_04294_),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_1 _09610_ (.A1(_02205_),
    .A2(_00072_),
    .B1(_04434_),
    .B2(_06534_),
    .X(_02246_));
 sky130_fd_sc_hd__nand4_1 _09611_ (.A(_02118_),
    .B(_02205_),
    .C(_04358_),
    .D(_00083_),
    .Y(_02247_));
 sky130_fd_sc_hd__a21bo_1 _09612_ (.A1(_02245_),
    .A2(_02246_),
    .B1_N(_02247_),
    .X(_02249_));
 sky130_fd_sc_hd__a21o_1 _09613_ (.A1(_02243_),
    .A2(_02244_),
    .B1(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__nand3_1 _09614_ (.A(_02243_),
    .B(_02244_),
    .C(_02249_),
    .Y(_02251_));
 sky130_fd_sc_hd__a21bo_1 _09615_ (.A1(_02242_),
    .A2(_02250_),
    .B1_N(_02251_),
    .X(_02252_));
 sky130_fd_sc_hd__and3_1 _09616_ (.A(_02238_),
    .B(_02239_),
    .C(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__xor2_1 _09617_ (.A(_02233_),
    .B(_02232_),
    .X(_02254_));
 sky130_fd_sc_hd__a21oi_1 _09618_ (.A1(_02238_),
    .A2(_02239_),
    .B1(_02252_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor3_2 _09619_ (.A(_02253_),
    .B(_02254_),
    .C(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__a21o_1 _09620_ (.A1(_02204_),
    .A2(_02207_),
    .B1(_02206_),
    .X(_02257_));
 sky130_fd_sc_hd__o211ai_2 _09621_ (.A1(_02253_),
    .A2(_02256_),
    .B1(_02208_),
    .C1(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__and3_1 _09622_ (.A(_02226_),
    .B(_02234_),
    .C(_02236_),
    .X(_02260_));
 sky130_fd_sc_hd__nor2_1 _09623_ (.A(_02237_),
    .B(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hd__a211o_1 _09624_ (.A1(_02208_),
    .A2(_02257_),
    .B1(_02253_),
    .C1(_02256_),
    .X(_02262_));
 sky130_fd_sc_hd__nand3_1 _09625_ (.A(_02258_),
    .B(_02261_),
    .C(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__o21a_1 _09626_ (.A1(_02211_),
    .A2(_02213_),
    .B1(_02212_),
    .X(_02264_));
 sky130_fd_sc_hd__a211o_1 _09627_ (.A1(_02258_),
    .A2(_02263_),
    .B1(_02214_),
    .C1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__o211ai_1 _09628_ (.A1(_02214_),
    .A2(_02264_),
    .B1(_02258_),
    .C1(_02263_),
    .Y(_02266_));
 sky130_fd_sc_hd__and3_1 _09629_ (.A(_02237_),
    .B(_02265_),
    .C(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__a21oi_1 _09630_ (.A1(_02265_),
    .A2(_02266_),
    .B1(_02237_),
    .Y(_02268_));
 sky130_fd_sc_hd__or2_1 _09631_ (.A(_02267_),
    .B(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__and4_1 _09632_ (.A(_06503_),
    .B(_06504_),
    .C(_00271_),
    .D(_04229_),
    .X(_02271_));
 sky130_fd_sc_hd__a22oi_2 _09633_ (.A1(_00162_),
    .A2(_00287_),
    .B1(_00267_),
    .B2(_00164_),
    .Y(_02272_));
 sky130_fd_sc_hd__and4bb_1 _09634_ (.A_N(_02272_),
    .B_N(_02271_),
    .C(_06475_),
    .D(_04111_),
    .X(_02273_));
 sky130_fd_sc_hd__nor2_1 _09635_ (.A(_02271_),
    .B(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _09636_ (.A(_02231_),
    .B(_02230_),
    .Y(_02275_));
 sky130_fd_sc_hd__xnor2_1 _09637_ (.A(_02228_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_1 _09638_ (.A(_02274_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_06560_),
    .B(_03873_),
    .Y(_02278_));
 sky130_fd_sc_hd__a22oi_1 _09640_ (.A1(_02229_),
    .A2(_06436_),
    .B1(_06446_),
    .B2(_02431_),
    .Y(_02279_));
 sky130_fd_sc_hd__and4_1 _09641_ (.A(_06520_),
    .B(_06516_),
    .C(net132),
    .D(_06430_),
    .X(_02280_));
 sky130_fd_sc_hd__o21ba_1 _09642_ (.A1(_02278_),
    .A2(_02279_),
    .B1_N(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__inv_2 _09643_ (.A(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__and2b_1 _09644_ (.A_N(_02274_),
    .B(_02276_),
    .X(_02283_));
 sky130_fd_sc_hd__a21oi_1 _09645_ (.A1(_02277_),
    .A2(_02282_),
    .B1(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__a22oi_1 _09646_ (.A1(_02669_),
    .A2(_03906_),
    .B1(_03993_),
    .B2(_02604_),
    .Y(_02285_));
 sky130_fd_sc_hd__or2_1 _09647_ (.A(_02169_),
    .B(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__nor2_1 _09648_ (.A(_02284_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(_02258_),
    .A2(_02262_),
    .B1(_02261_),
    .X(_02288_));
 sky130_fd_sc_hd__nand3_1 _09650_ (.A(_02251_),
    .B(_02242_),
    .C(_02250_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21o_1 _09651_ (.A1(_02251_),
    .A2(_02250_),
    .B1(_02242_),
    .X(_02290_));
 sky130_fd_sc_hd__o2bb2a_1 _09652_ (.A1_N(_06545_),
    .A2_N(_00303_),
    .B1(_02272_),
    .B2(_02271_),
    .X(_02292_));
 sky130_fd_sc_hd__nor2_1 _09653_ (.A(_02273_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand3_1 _09654_ (.A(_02247_),
    .B(_02245_),
    .C(_02246_),
    .Y(_02294_));
 sky130_fd_sc_hd__a22o_1 _09655_ (.A1(_02248_),
    .A2(_04305_),
    .B1(_02247_),
    .B2(_02246_),
    .X(_02295_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(_06488_),
    .B(_04229_),
    .Y(_02296_));
 sky130_fd_sc_hd__a22oi_2 _09657_ (.A1(_06463_),
    .A2(_00592_),
    .B1(_00072_),
    .B2(_06492_),
    .Y(_02297_));
 sky130_fd_sc_hd__and4_1 _09658_ (.A(_06469_),
    .B(_00150_),
    .C(net123),
    .D(_00089_),
    .X(_02298_));
 sky130_fd_sc_hd__o21bai_1 _09659_ (.A1(_02296_),
    .A2(_02297_),
    .B1_N(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__a21o_1 _09660_ (.A1(_02294_),
    .A2(_02295_),
    .B1(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__nand3_1 _09661_ (.A(_02294_),
    .B(_02295_),
    .C(_02299_),
    .Y(_02301_));
 sky130_fd_sc_hd__a21bo_1 _09662_ (.A1(_02293_),
    .A2(_02300_),
    .B1_N(_02301_),
    .X(_02303_));
 sky130_fd_sc_hd__nand3_2 _09663_ (.A(_02289_),
    .B(_02290_),
    .C(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__xnor2_1 _09664_ (.A(_02277_),
    .B(_02281_),
    .Y(_02305_));
 sky130_fd_sc_hd__a21o_1 _09665_ (.A1(_02289_),
    .A2(_02290_),
    .B1(_02303_),
    .X(_02306_));
 sky130_fd_sc_hd__nand3_2 _09666_ (.A(_02304_),
    .B(_02305_),
    .C(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__o21a_1 _09667_ (.A1(_02253_),
    .A2(_02255_),
    .B1(_02254_),
    .X(_02308_));
 sky130_fd_sc_hd__a211oi_4 _09668_ (.A1(_02304_),
    .A2(_02307_),
    .B1(_02256_),
    .C1(_02308_),
    .Y(_02309_));
 sky130_fd_sc_hd__xnor2_1 _09669_ (.A(_02284_),
    .B(_02286_),
    .Y(_02310_));
 sky130_fd_sc_hd__o211a_1 _09670_ (.A1(_02256_),
    .A2(_02308_),
    .B1(_02304_),
    .C1(_02307_),
    .X(_02311_));
 sky130_fd_sc_hd__nor3_1 _09671_ (.A(_02309_),
    .B(_02310_),
    .C(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__a211o_1 _09672_ (.A1(_02263_),
    .A2(_02288_),
    .B1(_02309_),
    .C1(_02312_),
    .X(_02314_));
 sky130_fd_sc_hd__o211ai_1 _09673_ (.A1(_02309_),
    .A2(_02312_),
    .B1(_02263_),
    .C1(_02288_),
    .Y(_02315_));
 sky130_fd_sc_hd__a21boi_1 _09674_ (.A1(_02287_),
    .A2(_02314_),
    .B1_N(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__or2_1 _09675_ (.A(_02269_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__and2b_1 _09676_ (.A_N(_02217_),
    .B(_02215_),
    .X(_02318_));
 sky130_fd_sc_hd__xnor2_1 _09677_ (.A(_02187_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__inv_2 _09678_ (.A(_02265_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _09679_ (.A(_02320_),
    .B(_02267_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_2 _09680_ (.A(_02319_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__or2_1 _09681_ (.A(_02317_),
    .B(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__or2_1 _09682_ (.A(_02219_),
    .B(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__a21boi_1 _09683_ (.A1(_02090_),
    .A2(_02163_),
    .B1_N(_02161_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21oi_1 _09684_ (.A1(_02916_),
    .A2(_03917_),
    .B1(_01918_),
    .Y(_02326_));
 sky130_fd_sc_hd__or2_1 _09685_ (.A(_01919_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__a21oi_1 _09686_ (.A1(_02153_),
    .A2(_02157_),
    .B1(_02327_),
    .Y(_02328_));
 sky130_fd_sc_hd__and3_1 _09687_ (.A(_02153_),
    .B(_02157_),
    .C(_02327_),
    .X(_02329_));
 sky130_fd_sc_hd__nor2_1 _09688_ (.A(_02328_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__a22o_1 _09689_ (.A1(_02014_),
    .A2(_02015_),
    .B1(_02016_),
    .B2(_01996_),
    .X(_02331_));
 sky130_fd_sc_hd__nand4_1 _09690_ (.A(_01996_),
    .B(_02014_),
    .C(_02015_),
    .D(_02016_),
    .Y(_02332_));
 sky130_fd_sc_hd__o211ai_1 _09691_ (.A1(_02147_),
    .A2(_02159_),
    .B1(_02331_),
    .C1(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__a211o_1 _09692_ (.A1(_02332_),
    .A2(_02331_),
    .B1(_02159_),
    .C1(_02147_),
    .X(_02335_));
 sky130_fd_sc_hd__and3_2 _09693_ (.A(_02330_),
    .B(_02333_),
    .C(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__a21oi_1 _09694_ (.A1(_02333_),
    .A2(_02335_),
    .B1(_02330_),
    .Y(_02337_));
 sky130_fd_sc_hd__or2_1 _09695_ (.A(_02336_),
    .B(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__xnor2_1 _09696_ (.A(_02325_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__xor2_2 _09697_ (.A(_02088_),
    .B(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__and2_1 _09698_ (.A(_02166_),
    .B(_02218_),
    .X(_02341_));
 sky130_fd_sc_hd__or2_1 _09699_ (.A(_02319_),
    .B(_02321_),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _09700_ (.A(_02219_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__or2_1 _09701_ (.A(_02341_),
    .B(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__xnor2_1 _09702_ (.A(_02340_),
    .B(_02344_),
    .Y(_02346_));
 sky130_fd_sc_hd__xnor2_2 _09703_ (.A(_02269_),
    .B(_02316_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand3_1 _09704_ (.A(_02301_),
    .B(_02293_),
    .C(_02300_),
    .Y(_02348_));
 sky130_fd_sc_hd__a21o_1 _09705_ (.A1(_02301_),
    .A2(_02300_),
    .B1(_02293_),
    .X(_02349_));
 sky130_fd_sc_hd__and2_1 _09706_ (.A(_06504_),
    .B(_04165_),
    .X(_02350_));
 sky130_fd_sc_hd__and2_1 _09707_ (.A(_06503_),
    .B(_04100_),
    .X(_02351_));
 sky130_fd_sc_hd__a22o_1 _09708_ (.A1(_02334_),
    .A2(_04100_),
    .B1(_00271_),
    .B2(_01332_),
    .X(_02352_));
 sky130_fd_sc_hd__a21bo_1 _09709_ (.A1(_02350_),
    .A2(_02351_),
    .B1_N(_02352_),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(_02377_),
    .B(_06443_),
    .Y(_02354_));
 sky130_fd_sc_hd__xor2_1 _09711_ (.A(_02353_),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__or3_1 _09712_ (.A(_02298_),
    .B(_02296_),
    .C(_02297_),
    .X(_02357_));
 sky130_fd_sc_hd__o21ai_1 _09713_ (.A1(_02298_),
    .A2(_02297_),
    .B1(_02296_),
    .Y(_02358_));
 sky130_fd_sc_hd__and2_1 _09714_ (.A(_06460_),
    .B(_04165_),
    .X(_02359_));
 sky130_fd_sc_hd__a22o_1 _09715_ (.A1(_00150_),
    .A2(net124),
    .B1(net123),
    .B2(_06469_),
    .X(_02360_));
 sky130_fd_sc_hd__nand4_1 _09716_ (.A(_06492_),
    .B(_06463_),
    .C(_00266_),
    .D(_00592_),
    .Y(_02361_));
 sky130_fd_sc_hd__a21bo_1 _09717_ (.A1(_02359_),
    .A2(_02360_),
    .B1_N(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__a21o_1 _09718_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__nand3_1 _09719_ (.A(_02357_),
    .B(_02358_),
    .C(_02362_),
    .Y(_02364_));
 sky130_fd_sc_hd__a21bo_1 _09720_ (.A1(_02355_),
    .A2(_02363_),
    .B1_N(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__and3_1 _09721_ (.A(_02348_),
    .B(_02349_),
    .C(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__a32o_1 _09722_ (.A1(_06545_),
    .A2(_04046_),
    .A3(_02352_),
    .B1(_02351_),
    .B2(_02350_),
    .X(_02367_));
 sky130_fd_sc_hd__nor2_1 _09723_ (.A(_02280_),
    .B(_02279_),
    .Y(_02368_));
 sky130_fd_sc_hd__xnor2_1 _09724_ (.A(_02278_),
    .B(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__xor2_1 _09725_ (.A(_02367_),
    .B(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__and4_1 _09726_ (.A(_02431_),
    .B(_02229_),
    .C(net115),
    .D(_06436_),
    .X(_02371_));
 sky130_fd_sc_hd__xnor2_1 _09727_ (.A(_02370_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__a21oi_1 _09728_ (.A1(_02348_),
    .A2(_02349_),
    .B1(_02365_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor3_2 _09729_ (.A(_02366_),
    .B(_02372_),
    .C(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__a21o_1 _09730_ (.A1(_02304_),
    .A2(_02306_),
    .B1(_02305_),
    .X(_02375_));
 sky130_fd_sc_hd__o211a_2 _09731_ (.A1(_02366_),
    .A2(_02374_),
    .B1(_02307_),
    .C1(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__and2_1 _09732_ (.A(_02367_),
    .B(_02369_),
    .X(_02378_));
 sky130_fd_sc_hd__and2_1 _09733_ (.A(_02370_),
    .B(_02371_),
    .X(_02379_));
 sky130_fd_sc_hd__o211a_1 _09734_ (.A1(_02378_),
    .A2(_02379_),
    .B1(_02604_),
    .C1(_03917_),
    .X(_02380_));
 sky130_fd_sc_hd__a211oi_1 _09735_ (.A1(_02604_),
    .A2(_03917_),
    .B1(_02378_),
    .C1(_02379_),
    .Y(_02381_));
 sky130_fd_sc_hd__or2_1 _09736_ (.A(_02380_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__a211oi_2 _09737_ (.A1(_02307_),
    .A2(_02375_),
    .B1(_02366_),
    .C1(_02374_),
    .Y(_02383_));
 sky130_fd_sc_hd__nor3_2 _09738_ (.A(_02376_),
    .B(_02382_),
    .C(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__or3_1 _09739_ (.A(_02309_),
    .B(_02310_),
    .C(_02311_),
    .X(_02385_));
 sky130_fd_sc_hd__o21ai_2 _09740_ (.A1(_02309_),
    .A2(_02311_),
    .B1(_02310_),
    .Y(_02386_));
 sky130_fd_sc_hd__o211ai_4 _09741_ (.A1(_02376_),
    .A2(_02384_),
    .B1(_02385_),
    .C1(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__a211o_1 _09742_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02376_),
    .C1(_02384_),
    .X(_02389_));
 sky130_fd_sc_hd__nand3_1 _09743_ (.A(_02380_),
    .B(_02387_),
    .C(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__and3_1 _09744_ (.A(_02287_),
    .B(_02315_),
    .C(_02314_),
    .X(_02391_));
 sky130_fd_sc_hd__a21oi_1 _09745_ (.A1(_02315_),
    .A2(_02314_),
    .B1(_02287_),
    .Y(_02392_));
 sky130_fd_sc_hd__a211oi_2 _09746_ (.A1(_02387_),
    .A2(_02390_),
    .B1(_02391_),
    .C1(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__inv_2 _09747_ (.A(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__or2_1 _09748_ (.A(_02347_),
    .B(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__and2_1 _09749_ (.A(_02342_),
    .B(_02323_),
    .X(_02396_));
 sky130_fd_sc_hd__xnor2_1 _09750_ (.A(_02219_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__nor3_1 _09751_ (.A(_02322_),
    .B(_02395_),
    .C(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__o21bai_1 _09752_ (.A1(_02324_),
    .A2(_02346_),
    .B1_N(_02398_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _09753_ (.A(_02322_),
    .B(_02395_),
    .Y(_02401_));
 sky130_fd_sc_hd__xor2_1 _09754_ (.A(_02401_),
    .B(_02397_),
    .X(_02402_));
 sky130_fd_sc_hd__o211a_1 _09755_ (.A1(_02391_),
    .A2(_02392_),
    .B1(_02387_),
    .C1(_02390_),
    .X(_02403_));
 sky130_fd_sc_hd__and3_1 _09756_ (.A(_02380_),
    .B(_02387_),
    .C(_02389_),
    .X(_02404_));
 sky130_fd_sc_hd__a21oi_1 _09757_ (.A1(_02387_),
    .A2(_02389_),
    .B1(_02380_),
    .Y(_02405_));
 sky130_fd_sc_hd__nor2_1 _09758_ (.A(_02404_),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3_1 _09759_ (.A(_02364_),
    .B(_02355_),
    .C(_02363_),
    .Y(_02407_));
 sky130_fd_sc_hd__a21o_1 _09760_ (.A1(_02364_),
    .A2(_02363_),
    .B1(_02355_),
    .X(_02408_));
 sky130_fd_sc_hd__and3_1 _09761_ (.A(_06479_),
    .B(net127),
    .C(net126),
    .X(_02409_));
 sky130_fd_sc_hd__a22o_1 _09762_ (.A1(_06480_),
    .A2(net127),
    .B1(net126),
    .B2(_06479_),
    .X(_02410_));
 sky130_fd_sc_hd__a21bo_1 _09763_ (.A1(_00162_),
    .A2(_02409_),
    .B1_N(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_06475_),
    .B(_03960_),
    .Y(_02412_));
 sky130_fd_sc_hd__xor2_1 _09765_ (.A(_02411_),
    .B(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__nand3_1 _09766_ (.A(_02361_),
    .B(_02359_),
    .C(_02360_),
    .Y(_02414_));
 sky130_fd_sc_hd__a22o_1 _09767_ (.A1(_02248_),
    .A2(_00287_),
    .B1(_02361_),
    .B2(_02360_),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_1 _09768_ (.A(net111),
    .B(net126),
    .Y(_02416_));
 sky130_fd_sc_hd__a22oi_2 _09769_ (.A1(_00150_),
    .A2(net125),
    .B1(_00266_),
    .B2(_06469_),
    .Y(_02417_));
 sky130_fd_sc_hd__and4_1 _09770_ (.A(_02096_),
    .B(net116),
    .C(net125),
    .D(net124),
    .X(_02418_));
 sky130_fd_sc_hd__o21bai_1 _09771_ (.A1(_02416_),
    .A2(_02417_),
    .B1_N(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21o_1 _09772_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02419_),
    .X(_02421_));
 sky130_fd_sc_hd__nand3_1 _09773_ (.A(_02414_),
    .B(_02415_),
    .C(_02419_),
    .Y(_02422_));
 sky130_fd_sc_hd__a21bo_1 _09774_ (.A1(_02413_),
    .A2(_02421_),
    .B1_N(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__nand3_2 _09775_ (.A(_02407_),
    .B(_02408_),
    .C(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__a22oi_1 _09776_ (.A1(_02229_),
    .A2(net115),
    .B1(_06437_),
    .B2(_02442_),
    .Y(_02425_));
 sky130_fd_sc_hd__or2_1 _09777_ (.A(_02371_),
    .B(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__and2_1 _09778_ (.A(_02345_),
    .B(_02409_),
    .X(_02427_));
 sky130_fd_sc_hd__a31o_1 _09779_ (.A1(_02388_),
    .A2(_03971_),
    .A3(_02410_),
    .B1(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__and2b_1 _09780_ (.A_N(_02426_),
    .B(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__and2b_1 _09781_ (.A_N(_02428_),
    .B(_02426_),
    .X(_02430_));
 sky130_fd_sc_hd__nor2_1 _09782_ (.A(_02429_),
    .B(_02430_),
    .Y(_02432_));
 sky130_fd_sc_hd__a21o_1 _09783_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02423_),
    .X(_02433_));
 sky130_fd_sc_hd__nand3_1 _09784_ (.A(_02424_),
    .B(_02432_),
    .C(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__o21a_1 _09785_ (.A1(_02366_),
    .A2(_02373_),
    .B1(_02372_),
    .X(_02435_));
 sky130_fd_sc_hd__a211oi_2 _09786_ (.A1(_02424_),
    .A2(_02434_),
    .B1(_02374_),
    .C1(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__o211a_1 _09787_ (.A1(_02374_),
    .A2(_02435_),
    .B1(_02424_),
    .C1(_02434_),
    .X(_02437_));
 sky130_fd_sc_hd__nor3b_2 _09788_ (.A(_02436_),
    .B(_02437_),
    .C_N(_02429_),
    .Y(_02438_));
 sky130_fd_sc_hd__or3_1 _09789_ (.A(_02376_),
    .B(_02382_),
    .C(_02383_),
    .X(_02439_));
 sky130_fd_sc_hd__o21ai_1 _09790_ (.A1(_02376_),
    .A2(_02383_),
    .B1(_02382_),
    .Y(_02440_));
 sky130_fd_sc_hd__o211a_1 _09791_ (.A1(_02436_),
    .A2(_02438_),
    .B1(_02439_),
    .C1(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__or4bb_1 _09792_ (.A(_02393_),
    .B(_02403_),
    .C_N(_02406_),
    .D_N(_02441_),
    .X(_02443_));
 sky130_fd_sc_hd__nor2_1 _09793_ (.A(_02347_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__o21ai_1 _09794_ (.A1(_02347_),
    .A2(_02394_),
    .B1(_02317_),
    .Y(_02445_));
 sky130_fd_sc_hd__xnor2_1 _09795_ (.A(_02322_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__or2_1 _09796_ (.A(_02444_),
    .B(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__inv_2 _09797_ (.A(_02406_),
    .Y(_02448_));
 sky130_fd_sc_hd__a211o_1 _09798_ (.A1(_02439_),
    .A2(_02440_),
    .B1(_02436_),
    .C1(_02438_),
    .X(_02449_));
 sky130_fd_sc_hd__nor2b_1 _09799_ (.A(_02441_),
    .B_N(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__nand3_1 _09800_ (.A(_02422_),
    .B(_02413_),
    .C(_02421_),
    .Y(_02451_));
 sky130_fd_sc_hd__a21o_1 _09801_ (.A1(_02422_),
    .A2(_02421_),
    .B1(_02413_),
    .X(_02452_));
 sky130_fd_sc_hd__a22oi_1 _09802_ (.A1(_06504_),
    .A2(net132),
    .B1(net127),
    .B2(_06503_),
    .Y(_02454_));
 sky130_fd_sc_hd__and4_1 _09803_ (.A(net110),
    .B(net109),
    .C(net132),
    .D(net127),
    .X(_02455_));
 sky130_fd_sc_hd__and4bb_1 _09804_ (.A_N(_02454_),
    .B_N(_02455_),
    .C(_06544_),
    .D(net115),
    .X(_02456_));
 sky130_fd_sc_hd__o2bb2a_1 _09805_ (.A1_N(_06544_),
    .A2_N(net115),
    .B1(_02454_),
    .B2(_02455_),
    .X(_02457_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_02456_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__or3_1 _09807_ (.A(_02418_),
    .B(_02416_),
    .C(_02417_),
    .X(_02459_));
 sky130_fd_sc_hd__o21ai_1 _09808_ (.A1(_02418_),
    .A2(_02417_),
    .B1(_02416_),
    .Y(_02460_));
 sky130_fd_sc_hd__a22o_1 _09809_ (.A1(_00150_),
    .A2(net126),
    .B1(net125),
    .B2(_06469_),
    .X(_02461_));
 sky130_fd_sc_hd__and4_1 _09810_ (.A(_06469_),
    .B(_00150_),
    .C(net126),
    .D(net125),
    .X(_02462_));
 sky130_fd_sc_hd__a31o_1 _09811_ (.A1(_02248_),
    .A2(_04035_),
    .A3(_02461_),
    .B1(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__a21o_1 _09812_ (.A1(_02459_),
    .A2(_02460_),
    .B1(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__and3_1 _09813_ (.A(_02459_),
    .B(_02460_),
    .C(_02463_),
    .X(_02465_));
 sky130_fd_sc_hd__a21o_1 _09814_ (.A1(_02458_),
    .A2(_02464_),
    .B1(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__and3_1 _09815_ (.A(_02451_),
    .B(_02452_),
    .C(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__inv_2 _09816_ (.A(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__o211a_1 _09817_ (.A1(_02455_),
    .A2(_02456_),
    .B1(_02442_),
    .C1(_03884_),
    .X(_02469_));
 sky130_fd_sc_hd__a211oi_1 _09818_ (.A1(_02442_),
    .A2(_03884_),
    .B1(_02455_),
    .C1(_02456_),
    .Y(_02470_));
 sky130_fd_sc_hd__or2_1 _09819_ (.A(_02469_),
    .B(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__a21oi_1 _09820_ (.A1(_02451_),
    .A2(_02452_),
    .B1(_02466_),
    .Y(_02472_));
 sky130_fd_sc_hd__or3_1 _09821_ (.A(_02467_),
    .B(_02471_),
    .C(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__and3_1 _09822_ (.A(_02424_),
    .B(_02432_),
    .C(_02433_),
    .X(_02475_));
 sky130_fd_sc_hd__a21oi_1 _09823_ (.A1(_02424_),
    .A2(_02433_),
    .B1(_02432_),
    .Y(_02476_));
 sky130_fd_sc_hd__a211o_1 _09824_ (.A1(_02468_),
    .A2(_02473_),
    .B1(_02475_),
    .C1(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__o211ai_1 _09825_ (.A1(_02475_),
    .A2(_02476_),
    .B1(_02468_),
    .C1(_02473_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand3_2 _09826_ (.A(_02469_),
    .B(_02477_),
    .C(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__o21ba_1 _09827_ (.A1(_02436_),
    .A2(_02437_),
    .B1_N(_02429_),
    .X(_02480_));
 sky130_fd_sc_hd__a211oi_2 _09828_ (.A1(_02477_),
    .A2(_02479_),
    .B1(_02438_),
    .C1(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(_02450_),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__a2bb2o_1 _09830_ (.A1_N(_02393_),
    .A2_N(_02403_),
    .B1(_02406_),
    .B2(_02441_),
    .X(_02483_));
 sky130_fd_sc_hd__or4bb_1 _09831_ (.A(_02448_),
    .B(_02482_),
    .C_N(_02483_),
    .D_N(_02443_),
    .X(_02484_));
 sky130_fd_sc_hd__a2bb2o_1 _09832_ (.A1_N(_02448_),
    .A2_N(_02482_),
    .B1(_02483_),
    .B2(_02443_),
    .X(_02486_));
 sky130_fd_sc_hd__a21o_1 _09833_ (.A1(_02449_),
    .A2(_02481_),
    .B1(_02441_),
    .X(_02487_));
 sky130_fd_sc_hd__or3_1 _09834_ (.A(_02404_),
    .B(_02405_),
    .C(_02487_),
    .X(_02488_));
 sky130_fd_sc_hd__o21ai_1 _09835_ (.A1(_02404_),
    .A2(_02405_),
    .B1(_02487_),
    .Y(_02489_));
 sky130_fd_sc_hd__a211o_1 _09836_ (.A1(_02477_),
    .A2(_02479_),
    .B1(_02438_),
    .C1(_02480_),
    .X(_02490_));
 sky130_fd_sc_hd__o211ai_1 _09837_ (.A1(_02438_),
    .A2(_02480_),
    .B1(_02477_),
    .C1(_02479_),
    .Y(_02491_));
 sky130_fd_sc_hd__a21o_1 _09838_ (.A1(_02477_),
    .A2(_02478_),
    .B1(_02469_),
    .X(_02492_));
 sky130_fd_sc_hd__and4_1 _09839_ (.A(_06492_),
    .B(_06463_),
    .C(net127),
    .D(_04100_),
    .X(_02493_));
 sky130_fd_sc_hd__a22oi_2 _09840_ (.A1(_02205_),
    .A2(_06430_),
    .B1(_06431_),
    .B2(_06534_),
    .Y(_02494_));
 sky130_fd_sc_hd__and4bb_1 _09841_ (.A_N(_02493_),
    .B_N(_02494_),
    .C(_02248_),
    .D(_03960_),
    .X(_02495_));
 sky130_fd_sc_hd__nor2_1 _09842_ (.A(_02493_),
    .B(_02495_),
    .Y(_02497_));
 sky130_fd_sc_hd__nand2_1 _09843_ (.A(_02248_),
    .B(_06446_),
    .Y(_02498_));
 sky130_fd_sc_hd__and2b_1 _09844_ (.A_N(_02462_),
    .B(_02461_),
    .X(_02499_));
 sky130_fd_sc_hd__xnor2_1 _09845_ (.A(_02498_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__or2b_1 _09846_ (.A(_02497_),
    .B_N(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__a22o_1 _09847_ (.A1(_02345_),
    .A2(_03873_),
    .B1(_03971_),
    .B2(_02302_),
    .X(_02502_));
 sky130_fd_sc_hd__and4_1 _09848_ (.A(_02302_),
    .B(_02345_),
    .C(net115),
    .D(_06436_),
    .X(_02503_));
 sky130_fd_sc_hd__inv_2 _09849_ (.A(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_02502_),
    .B(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__xnor2_1 _09851_ (.A(_02500_),
    .B(_02497_),
    .Y(_02506_));
 sky130_fd_sc_hd__or2b_1 _09852_ (.A(_02505_),
    .B_N(_02506_),
    .X(_02508_));
 sky130_fd_sc_hd__and2b_1 _09853_ (.A_N(_02465_),
    .B(_02464_),
    .X(_02509_));
 sky130_fd_sc_hd__xnor2_1 _09854_ (.A(_02458_),
    .B(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__a21o_1 _09855_ (.A1(_02501_),
    .A2(_02508_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__and3_1 _09856_ (.A(_02510_),
    .B(_02501_),
    .C(_02508_),
    .X(_02512_));
 sky130_fd_sc_hd__or3b_1 _09857_ (.A(_02512_),
    .B(_02504_),
    .C_N(_02511_),
    .X(_02513_));
 sky130_fd_sc_hd__o21ai_1 _09858_ (.A1(_02467_),
    .A2(_02472_),
    .B1(_02471_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_1 _09859_ (.A(_02473_),
    .B(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__a21oi_1 _09860_ (.A1(_02511_),
    .A2(_02513_),
    .B1(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__and3_1 _09861_ (.A(_02479_),
    .B(_02492_),
    .C(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__and3_1 _09862_ (.A(_02490_),
    .B(_02491_),
    .C(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(_02450_),
    .B(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a21oi_1 _09864_ (.A1(_02488_),
    .A2(_02489_),
    .B1(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21o_1 _09865_ (.A1(_02484_),
    .A2(_02486_),
    .B1(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__a21o_1 _09866_ (.A1(_02488_),
    .A2(_02489_),
    .B1(_02519_),
    .X(_02522_));
 sky130_fd_sc_hd__nand3_1 _09867_ (.A(_02519_),
    .B(_02488_),
    .C(_02489_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(_02479_),
    .B(_02492_),
    .Y(_02524_));
 sky130_fd_sc_hd__a21oi_1 _09869_ (.A1(_02490_),
    .A2(_02491_),
    .B1(_02517_),
    .Y(_02525_));
 sky130_fd_sc_hd__and3_1 _09870_ (.A(_02515_),
    .B(_02511_),
    .C(_02513_),
    .X(_02526_));
 sky130_fd_sc_hd__a21oi_1 _09871_ (.A1(_02501_),
    .A2(_02508_),
    .B1(_02510_),
    .Y(_02527_));
 sky130_fd_sc_hd__or2_1 _09872_ (.A(_02527_),
    .B(_02512_),
    .X(_02529_));
 sky130_fd_sc_hd__xnor2_1 _09873_ (.A(_02503_),
    .B(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__and4_1 _09874_ (.A(_02118_),
    .B(_02216_),
    .C(_06437_),
    .D(_04046_),
    .X(_02531_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_02216_),
    .B(_06437_),
    .Y(_02532_));
 sky130_fd_sc_hd__a21boi_1 _09876_ (.A1(_02118_),
    .A2(_04057_),
    .B1_N(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__nor2_1 _09877_ (.A(_02531_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__and3_1 _09878_ (.A(_02259_),
    .B(_03895_),
    .C(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__o2bb2a_1 _09879_ (.A1_N(_02259_),
    .A2_N(_03982_),
    .B1(_02493_),
    .B2(_02494_),
    .X(_02536_));
 sky130_fd_sc_hd__nor2_1 _09880_ (.A(_02495_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__o21a_1 _09881_ (.A1(_02531_),
    .A2(_02535_),
    .B1(_02537_),
    .X(_02538_));
 sky130_fd_sc_hd__nor3_1 _09882_ (.A(_02537_),
    .B(_02531_),
    .C(_02535_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor2_1 _09883_ (.A(_02538_),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__and3_1 _09884_ (.A(_02302_),
    .B(_03917_),
    .C(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__xnor2_1 _09885_ (.A(_02505_),
    .B(_02506_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21a_1 _09886_ (.A1(_02538_),
    .A2(_02542_),
    .B1(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__or4bb_1 _09887_ (.A(_02516_),
    .B(_02526_),
    .C_N(_02530_),
    .D_N(_02544_),
    .X(_02545_));
 sky130_fd_sc_hd__or4_2 _09888_ (.A(_02524_),
    .B(_02518_),
    .C(_02525_),
    .D(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__a21oi_1 _09889_ (.A1(_02491_),
    .A2(_02517_),
    .B1(_02481_),
    .Y(_02547_));
 sky130_fd_sc_hd__xnor2_1 _09890_ (.A(_02450_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__and2b_1 _09891_ (.A_N(_02546_),
    .B(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__a21o_1 _09892_ (.A1(_02522_),
    .A2(_02523_),
    .B1(_02549_),
    .X(_02551_));
 sky130_fd_sc_hd__nand2_1 _09893_ (.A(_02530_),
    .B(_02544_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21ai_1 _09894_ (.A1(_02516_),
    .A2(_02526_),
    .B1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor3_1 _09895_ (.A(_02543_),
    .B(_02538_),
    .C(_02542_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _09896_ (.A(_02302_),
    .B(_03928_),
    .Y(_02555_));
 sky130_fd_sc_hd__xnor2_1 _09897_ (.A(_02555_),
    .B(_02541_),
    .Y(_02556_));
 sky130_fd_sc_hd__a21o_1 _09898_ (.A1(_02259_),
    .A2(_03917_),
    .B1(_02534_),
    .X(_02557_));
 sky130_fd_sc_hd__and2b_1 _09899_ (.A_N(_02535_),
    .B(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_2 _09900_ (.A(_02118_),
    .B(_03895_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _09901_ (.A(_02532_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__and2_1 _09902_ (.A(_02558_),
    .B(_02560_),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_1 _09903_ (.A(_02556_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor3_1 _09904_ (.A(_02544_),
    .B(_02554_),
    .C(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__and2_1 _09905_ (.A(_02530_),
    .B(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__nand3_1 _09906_ (.A(_02545_),
    .B(_02553_),
    .C(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hd__or2b_1 _09907_ (.A(_02516_),
    .B_N(_02545_),
    .X(_02567_));
 sky130_fd_sc_hd__xor2_1 _09908_ (.A(_02524_),
    .B(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__o22ai_1 _09909_ (.A1(_02518_),
    .A2(_02525_),
    .B1(_02545_),
    .B2(_02524_),
    .Y(_02569_));
 sky130_fd_sc_hd__and4bb_1 _09910_ (.A_N(_02566_),
    .B_N(_02568_),
    .C(_02546_),
    .D(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__and2_1 _09911_ (.A(_02548_),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__and3_1 _09912_ (.A(_02522_),
    .B(_02523_),
    .C(_02549_),
    .X(_02572_));
 sky130_fd_sc_hd__a21o_1 _09913_ (.A1(_02551_),
    .A2(_02571_),
    .B1(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__and3_1 _09914_ (.A(_02484_),
    .B(_02486_),
    .C(_02520_),
    .X(_02574_));
 sky130_fd_sc_hd__a21o_1 _09915_ (.A1(_02521_),
    .A2(_02573_),
    .B1(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__and3_1 _09916_ (.A(_02347_),
    .B(_02394_),
    .C(_02443_),
    .X(_02576_));
 sky130_fd_sc_hd__a21oi_1 _09917_ (.A1(_02394_),
    .A2(_02443_),
    .B1(_02347_),
    .Y(_02577_));
 sky130_fd_sc_hd__or2_1 _09918_ (.A(_02576_),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__xor2_1 _09919_ (.A(_02484_),
    .B(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__and2_1 _09920_ (.A(_02444_),
    .B(_02446_),
    .X(_02580_));
 sky130_fd_sc_hd__nor2_1 _09921_ (.A(_02484_),
    .B(_02578_),
    .Y(_02581_));
 sky130_fd_sc_hd__a211o_1 _09922_ (.A1(_02575_),
    .A2(_02579_),
    .B1(_02580_),
    .C1(_02581_),
    .X(_02583_));
 sky130_fd_sc_hd__and3b_2 _09923_ (.A_N(_02402_),
    .B(_02447_),
    .C(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__or2b_1 _09924_ (.A(_01959_),
    .B_N(_01964_),
    .X(_02585_));
 sky130_fd_sc_hd__o211a_1 _09925_ (.A1(_02147_),
    .A2(_02159_),
    .B1(_02331_),
    .C1(_02332_),
    .X(_02586_));
 sky130_fd_sc_hd__a21o_1 _09926_ (.A1(_02021_),
    .A2(_02027_),
    .B1(_02026_),
    .X(_02587_));
 sky130_fd_sc_hd__o211ai_4 _09927_ (.A1(_02586_),
    .A2(_02336_),
    .B1(_02587_),
    .C1(_02028_),
    .Y(_02588_));
 sky130_fd_sc_hd__a211o_1 _09928_ (.A1(_02028_),
    .A2(_02587_),
    .B1(_02336_),
    .C1(_02586_),
    .X(_02589_));
 sky130_fd_sc_hd__nand3_1 _09929_ (.A(_02328_),
    .B(_02588_),
    .C(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__o21ba_1 _09930_ (.A1(_02032_),
    .A2(_02033_),
    .B1_N(_02024_),
    .X(_02591_));
 sky130_fd_sc_hd__a211oi_2 _09931_ (.A1(_02588_),
    .A2(_02590_),
    .B1(_02591_),
    .C1(_02034_),
    .Y(_02592_));
 sky130_fd_sc_hd__a211o_1 _09932_ (.A1(_02035_),
    .A2(_02036_),
    .B1(_02032_),
    .C1(_02034_),
    .X(_02594_));
 sky130_fd_sc_hd__a21oi_1 _09933_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02037_),
    .Y(_02595_));
 sky130_fd_sc_hd__xnor2_1 _09934_ (.A(_02585_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__or2b_1 _09935_ (.A(_02037_),
    .B_N(_02594_),
    .X(_02597_));
 sky130_fd_sc_hd__or3_1 _09936_ (.A(_02325_),
    .B(_02336_),
    .C(_02337_),
    .X(_02598_));
 sky130_fd_sc_hd__o21a_1 _09937_ (.A1(_02336_),
    .A2(_02337_),
    .B1(_02325_),
    .X(_02599_));
 sky130_fd_sc_hd__or3b_1 _09938_ (.A(_02599_),
    .B(_02088_),
    .C_N(_02598_),
    .X(_02600_));
 sky130_fd_sc_hd__and3_1 _09939_ (.A(_02328_),
    .B(_02588_),
    .C(_02589_),
    .X(_02601_));
 sky130_fd_sc_hd__a21oi_1 _09940_ (.A1(_02588_),
    .A2(_02589_),
    .B1(_02328_),
    .Y(_02602_));
 sky130_fd_sc_hd__a211o_1 _09941_ (.A1(_02598_),
    .A2(_02600_),
    .B1(_02601_),
    .C1(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__o211a_1 _09942_ (.A1(_02034_),
    .A2(_02591_),
    .B1(_02590_),
    .C1(_02588_),
    .X(_02605_));
 sky130_fd_sc_hd__o21ba_1 _09943_ (.A1(_02603_),
    .A2(_02605_),
    .B1_N(_02592_),
    .X(_02606_));
 sky130_fd_sc_hd__xnor2_1 _09944_ (.A(_02597_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__or2_1 _09945_ (.A(_02596_),
    .B(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__or2_2 _09946_ (.A(_02592_),
    .B(_02605_),
    .X(_02609_));
 sky130_fd_sc_hd__o211ai_2 _09947_ (.A1(_02601_),
    .A2(_02602_),
    .B1(_02598_),
    .C1(_02600_),
    .Y(_02610_));
 sky130_fd_sc_hd__a211oi_1 _09948_ (.A1(_02598_),
    .A2(_02600_),
    .B1(_02601_),
    .C1(_02602_),
    .Y(_02611_));
 sky130_fd_sc_hd__a31o_1 _09949_ (.A1(_02341_),
    .A2(_02340_),
    .A3(_02610_),
    .B1(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__xnor2_2 _09950_ (.A(_02609_),
    .B(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand4_1 _09951_ (.A(_02341_),
    .B(_02340_),
    .C(_02603_),
    .D(_02610_),
    .Y(_02614_));
 sky130_fd_sc_hd__a22o_1 _09952_ (.A1(_02341_),
    .A2(_02340_),
    .B1(_02603_),
    .B2(_02610_),
    .X(_02616_));
 sky130_fd_sc_hd__and2_1 _09953_ (.A(_02614_),
    .B(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__and2_1 _09954_ (.A(_02340_),
    .B(_02343_),
    .X(_02618_));
 sky130_fd_sc_hd__xor2_2 _09955_ (.A(_02617_),
    .B(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__and3b_1 _09956_ (.A_N(_02608_),
    .B(_02613_),
    .C(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_02324_),
    .B(_02346_),
    .Y(_02621_));
 sky130_fd_sc_hd__o211a_1 _09958_ (.A1(_02400_),
    .A2(_02584_),
    .B1(_02620_),
    .C1(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__nor2_1 _09959_ (.A(_02614_),
    .B(_02609_),
    .Y(_02623_));
 sky130_fd_sc_hd__a31oi_1 _09960_ (.A1(_02617_),
    .A2(_02618_),
    .A3(_02613_),
    .B1(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__clkinv_2 _09961_ (.A(_02592_),
    .Y(_02625_));
 sky130_fd_sc_hd__or3_1 _09962_ (.A(_02585_),
    .B(_02625_),
    .C(_02597_),
    .X(_02627_));
 sky130_fd_sc_hd__or3_1 _09963_ (.A(_02603_),
    .B(_02597_),
    .C(_02609_),
    .X(_02628_));
 sky130_fd_sc_hd__or2_1 _09964_ (.A(_02596_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__o211ai_1 _09965_ (.A1(_02608_),
    .A2(_02624_),
    .B1(_02627_),
    .C1(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__and2_1 _09966_ (.A(_02041_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__nand3b_2 _09967_ (.A_N(_01676_),
    .B(_01767_),
    .C(_01844_),
    .Y(_02632_));
 sky130_fd_sc_hd__inv_2 _09968_ (.A(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__or2_1 _09969_ (.A(_01676_),
    .B(_01845_),
    .X(_02634_));
 sky130_fd_sc_hd__o211ai_2 _09970_ (.A1(_01848_),
    .A2(_01849_),
    .B1(_01878_),
    .C1(_01879_),
    .Y(_02635_));
 sky130_fd_sc_hd__a211o_1 _09971_ (.A1(_01878_),
    .A2(_01879_),
    .B1(_01848_),
    .C1(_01849_),
    .X(_02636_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(_02635_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_02634_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__and3_1 _09974_ (.A(_01767_),
    .B(_01959_),
    .C(_01963_),
    .X(_02639_));
 sky130_fd_sc_hd__or4bb_1 _09975_ (.A(_01844_),
    .B(_02585_),
    .C_N(_02037_),
    .D_N(_01960_),
    .X(_02640_));
 sky130_fd_sc_hd__nor2_1 _09976_ (.A(_01962_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__o211a_1 _09977_ (.A1(_02639_),
    .A2(_02641_),
    .B1(_01847_),
    .C1(_01881_),
    .X(_02642_));
 sky130_fd_sc_hd__nor2_1 _09978_ (.A(_02634_),
    .B(_02637_),
    .Y(_02643_));
 sky130_fd_sc_hd__a211o_1 _09979_ (.A1(_02633_),
    .A2(_02638_),
    .B1(_02642_),
    .C1(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__a211o_4 _09980_ (.A1(_02041_),
    .A2(_02622_),
    .B1(_02631_),
    .C1(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__o211ai_2 _09981_ (.A1(_01631_),
    .A2(_01852_),
    .B1(_01853_),
    .C1(_01854_),
    .Y(_02646_));
 sky130_fd_sc_hd__a22oi_4 _09982_ (.A1(_01304_),
    .A2(_01305_),
    .B1(_01306_),
    .B2(_01307_),
    .Y(_02648_));
 sky130_fd_sc_hd__and4_1 _09983_ (.A(_01304_),
    .B(_01305_),
    .C(_01306_),
    .D(_01307_),
    .X(_02649_));
 sky130_fd_sc_hd__a211oi_4 _09984_ (.A1(_02646_),
    .A2(_01865_),
    .B1(_02648_),
    .C1(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__or2_1 _09985_ (.A(_01860_),
    .B(_01862_),
    .X(_02651_));
 sky130_fd_sc_hd__xnor2_1 _09986_ (.A(_01871_),
    .B(_01213_),
    .Y(_02652_));
 sky130_fd_sc_hd__xnor2_1 _09987_ (.A(_02651_),
    .B(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__o211a_1 _09988_ (.A1(_02649_),
    .A2(_02648_),
    .B1(_01865_),
    .C1(_02646_),
    .X(_02654_));
 sky130_fd_sc_hd__nor3_1 _09989_ (.A(_02650_),
    .B(_02653_),
    .C(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__o21ai_1 _09990_ (.A1(_01311_),
    .A2(_01312_),
    .B1(_01313_),
    .Y(_02656_));
 sky130_fd_sc_hd__or3_1 _09991_ (.A(_01311_),
    .B(_01312_),
    .C(_01313_),
    .X(_02657_));
 sky130_fd_sc_hd__o211ai_2 _09992_ (.A1(_02650_),
    .A2(_02655_),
    .B1(_02656_),
    .C1(_02657_),
    .Y(_02659_));
 sky130_fd_sc_hd__and2_1 _09993_ (.A(_02651_),
    .B(_02652_),
    .X(_02660_));
 sky130_fd_sc_hd__a211o_1 _09994_ (.A1(_02657_),
    .A2(_02656_),
    .B1(_02655_),
    .C1(_02650_),
    .X(_02661_));
 sky130_fd_sc_hd__nand3_1 _09995_ (.A(_02660_),
    .B(_02659_),
    .C(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a21oi_1 _09996_ (.A1(_01316_),
    .A2(_01315_),
    .B1(_01275_),
    .Y(_02663_));
 sky130_fd_sc_hd__and3_1 _09997_ (.A(_01316_),
    .B(_01275_),
    .C(_01315_),
    .X(_02664_));
 sky130_fd_sc_hd__a211o_2 _09998_ (.A1(_02659_),
    .A2(_02662_),
    .B1(_02663_),
    .C1(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__o211ai_1 _09999_ (.A1(_02664_),
    .A2(_02663_),
    .B1(_02662_),
    .C1(_02659_),
    .Y(_02666_));
 sky130_fd_sc_hd__nor3_1 _10000_ (.A(_01866_),
    .B(_01867_),
    .C(_01873_),
    .Y(_02667_));
 sky130_fd_sc_hd__o21ai_1 _10001_ (.A1(_02650_),
    .A2(_02654_),
    .B1(_02653_),
    .Y(_02668_));
 sky130_fd_sc_hd__or3_1 _10002_ (.A(_02650_),
    .B(_02653_),
    .C(_02654_),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_1 _10003_ (.A1(_01866_),
    .A2(_02667_),
    .B1(_02668_),
    .C1(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__nand2_1 _10004_ (.A(_01868_),
    .B(_01872_),
    .Y(_02672_));
 sky130_fd_sc_hd__a211oi_1 _10005_ (.A1(_02670_),
    .A2(_02668_),
    .B1(_02667_),
    .C1(_01866_),
    .Y(_02673_));
 sky130_fd_sc_hd__nor3_2 _10006_ (.A(_02672_),
    .B(_02671_),
    .C(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21o_1 _10007_ (.A1(_02659_),
    .A2(_02661_),
    .B1(_02660_),
    .X(_02675_));
 sky130_fd_sc_hd__o211a_1 _10008_ (.A1(_02671_),
    .A2(_02674_),
    .B1(_02675_),
    .C1(_02662_),
    .X(_02676_));
 sky130_fd_sc_hd__nand3_1 _10009_ (.A(_02665_),
    .B(_02666_),
    .C(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__a21o_1 _10010_ (.A1(_02665_),
    .A2(_02666_),
    .B1(_02676_),
    .X(_02678_));
 sky130_fd_sc_hd__and2_1 _10011_ (.A(_02677_),
    .B(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__a21oi_1 _10012_ (.A1(_01202_),
    .A2(_01318_),
    .B1(_01317_),
    .Y(_02681_));
 sky130_fd_sc_hd__nor2_2 _10013_ (.A(_01319_),
    .B(_02681_),
    .Y(_02682_));
 sky130_fd_sc_hd__xnor2_4 _10014_ (.A(_02665_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__o21a_1 _10015_ (.A1(_02671_),
    .A2(_02673_),
    .B1(_02672_),
    .X(_02684_));
 sky130_fd_sc_hd__a211oi_2 _10016_ (.A1(_01876_),
    .A2(_01878_),
    .B1(_02684_),
    .C1(_02674_),
    .Y(_02685_));
 sky130_fd_sc_hd__o211a_1 _10017_ (.A1(_02674_),
    .A2(_02684_),
    .B1(_01878_),
    .C1(_01876_),
    .X(_02686_));
 sky130_fd_sc_hd__nor3_1 _10018_ (.A(_02635_),
    .B(_02685_),
    .C(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__o21a_1 _10019_ (.A1(_02685_),
    .A2(_02686_),
    .B1(_02635_),
    .X(_02688_));
 sky130_fd_sc_hd__a211oi_1 _10020_ (.A1(_02662_),
    .A2(_02675_),
    .B1(_02674_),
    .C1(_02671_),
    .Y(_02689_));
 sky130_fd_sc_hd__nor2_1 _10021_ (.A(_02676_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__xnor2_1 _10022_ (.A(_02685_),
    .B(_02690_),
    .Y(_02692_));
 sky130_fd_sc_hd__nor3_1 _10023_ (.A(_02687_),
    .B(_02688_),
    .C(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__and3_1 _10024_ (.A(_02679_),
    .B(_02683_),
    .C(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__and2_1 _10025_ (.A(_00817_),
    .B(_00818_),
    .X(_02695_));
 sky130_fd_sc_hd__o21ai_1 _10026_ (.A1(_01328_),
    .A2(_01329_),
    .B1(_00954_),
    .Y(_02696_));
 sky130_fd_sc_hd__o21a_1 _10027_ (.A1(_02685_),
    .A2(_02687_),
    .B1(_02690_),
    .X(_02697_));
 sky130_fd_sc_hd__nand2_1 _10028_ (.A(_02665_),
    .B(_02677_),
    .Y(_02698_));
 sky130_fd_sc_hd__a32o_2 _10029_ (.A1(_02679_),
    .A2(_02683_),
    .A3(_02697_),
    .B1(_02698_),
    .B2(_02682_),
    .X(_02699_));
 sky130_fd_sc_hd__a21oi_1 _10030_ (.A1(_01200_),
    .A2(_01320_),
    .B1(_01326_),
    .Y(_02700_));
 sky130_fd_sc_hd__o211a_1 _10031_ (.A1(_00955_),
    .A2(_00956_),
    .B1(_02700_),
    .C1(_01330_),
    .X(_02701_));
 sky130_fd_sc_hd__a221o_1 _10032_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02699_),
    .B2(_01331_),
    .C1(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__a31o_4 _10033_ (.A1(_01331_),
    .A2(_02645_),
    .A3(_02694_),
    .B1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__xor2_2 _10034_ (.A(_00816_),
    .B(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__clkbuf_4 _10035_ (.A(net2),
    .X(_02705_));
 sky130_fd_sc_hd__or2b_1 _10036_ (.A(net4),
    .B_N(net3),
    .X(_02706_));
 sky130_fd_sc_hd__nor2_2 _10037_ (.A(_02064_),
    .B(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nand2_1 _10038_ (.A(_02705_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__nand2_1 _10039_ (.A(_02705_),
    .B(_02020_),
    .Y(_02709_));
 sky130_fd_sc_hd__or3b_1 _10040_ (.A(_06023_),
    .B(_02709_),
    .C_N(_02064_),
    .X(_02710_));
 sky130_fd_sc_hd__buf_2 _10041_ (.A(_02710_),
    .X(_02711_));
 sky130_fd_sc_hd__nand3_4 _10042_ (.A(_02020_),
    .B(_06023_),
    .C(_02075_),
    .Y(_02713_));
 sky130_fd_sc_hd__or2b_1 _10043_ (.A(_02118_),
    .B_N(_03917_),
    .X(_02714_));
 sky130_fd_sc_hd__nand2b_2 _10044_ (.A_N(_03906_),
    .B(_02118_),
    .Y(_02715_));
 sky130_fd_sc_hd__a32o_1 _10045_ (.A1(_02708_),
    .A2(_02711_),
    .A3(_02713_),
    .B1(_02714_),
    .B2(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__and3b_1 _10046_ (.A_N(_06023_),
    .B(_02075_),
    .C(_02020_),
    .X(_02717_));
 sky130_fd_sc_hd__clkbuf_4 _10047_ (.A(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__buf_4 _10048_ (.A(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__or2_2 _10049_ (.A(_02064_),
    .B(_02706_),
    .X(_02720_));
 sky130_fd_sc_hd__nor2_4 _10050_ (.A(_02705_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__clkbuf_4 _10051_ (.A(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__clkbuf_4 _10052_ (.A(_02722_),
    .X(_02724_));
 sky130_fd_sc_hd__o21a_1 _10053_ (.A1(_02118_),
    .A2(_03928_),
    .B1(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__or3_2 _10054_ (.A(_02064_),
    .B(net3),
    .C(_02709_),
    .X(_02726_));
 sky130_fd_sc_hd__clkbuf_4 _10055_ (.A(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_2 _10056_ (.A(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__and2_1 _10057_ (.A(net2),
    .B(net1),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_1 _10058_ (.A1(_02075_),
    .A2(_02729_),
    .B1(_02031_),
    .X(_02730_));
 sky130_fd_sc_hd__buf_2 _10059_ (.A(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__clkbuf_4 _10060_ (.A(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__a2bb2o_1 _10061_ (.A1_N(_03928_),
    .A2_N(_02728_),
    .B1(_02732_),
    .B2(\AuI.result[0] ),
    .X(_02733_));
 sky130_fd_sc_hd__a211o_1 _10062_ (.A1(_04004_),
    .A2(_02719_),
    .B1(_02725_),
    .C1(_02733_),
    .X(_02735_));
 sky130_fd_sc_hd__and3_2 _10063_ (.A(_02129_),
    .B(_02064_),
    .C(_02031_),
    .X(_02736_));
 sky130_fd_sc_hd__clkbuf_4 _10064_ (.A(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__clkbuf_4 _10065_ (.A(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_4 _10066_ (.A(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__and4b_1 _10067_ (.A_N(_02064_),
    .B(_02020_),
    .C(_06023_),
    .D(_02705_),
    .X(_02740_));
 sky130_fd_sc_hd__buf_6 _10068_ (.A(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__and3b_1 _10069_ (.A_N(_02706_),
    .B(_02129_),
    .C(_02064_),
    .X(_02742_));
 sky130_fd_sc_hd__buf_2 _10070_ (.A(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__buf_2 _10071_ (.A(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__clkbuf_4 _10072_ (.A(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__o21ba_1 _10073_ (.A1(_02741_),
    .A2(_02745_),
    .B1_N(_02559_),
    .X(_02746_));
 sky130_fd_sc_hd__a221o_1 _10074_ (.A1(\MuI.result[0] ),
    .A2(_02739_),
    .B1(_06056_),
    .B2(\FuI.Integer[0] ),
    .C1(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__nor2_1 _10075_ (.A(_02735_),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__o211ai_4 _10076_ (.A1(_06428_),
    .A2(_02704_),
    .B1(_02716_),
    .C1(_02748_),
    .Y(net69));
 sky130_fd_sc_hd__and3_1 _10077_ (.A(_02020_),
    .B(_06023_),
    .C(_02075_),
    .X(_02749_));
 sky130_fd_sc_hd__clkbuf_4 _10078_ (.A(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__buf_6 _10079_ (.A(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__buf_4 _10080_ (.A(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__xnor2_4 _10081_ (.A(_02216_),
    .B(_03982_),
    .Y(_02753_));
 sky130_fd_sc_hd__xnor2_1 _10082_ (.A(_02715_),
    .B(_02753_),
    .Y(_02755_));
 sky130_fd_sc_hd__or2_1 _10083_ (.A(_02442_),
    .B(_04327_),
    .X(_02756_));
 sky130_fd_sc_hd__nand2_2 _10084_ (.A(_01988_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__and2b_1 _10085_ (.A_N(_04251_),
    .B(_02388_),
    .X(_02758_));
 sky130_fd_sc_hd__and2b_1 _10086_ (.A_N(_02388_),
    .B(_04262_),
    .X(_02759_));
 sky130_fd_sc_hd__nor2_2 _10087_ (.A(_02758_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__and2b_1 _10088_ (.A_N(_02345_),
    .B(_04186_),
    .X(_02761_));
 sky130_fd_sc_hd__and2b_1 _10089_ (.A_N(_04186_),
    .B(_02345_),
    .X(_02762_));
 sky130_fd_sc_hd__or2_1 _10090_ (.A(_02761_),
    .B(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__buf_2 _10091_ (.A(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__inv_2 _10092_ (.A(_02764_),
    .Y(_02766_));
 sky130_fd_sc_hd__xnor2_4 _10093_ (.A(_02259_),
    .B(_04057_),
    .Y(_02767_));
 sky130_fd_sc_hd__xnor2_1 _10094_ (.A(_02302_),
    .B(_04122_),
    .Y(_02768_));
 sky130_fd_sc_hd__and2_1 _10095_ (.A(_02767_),
    .B(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__and3_1 _10096_ (.A(_02715_),
    .B(_02714_),
    .C(_02753_),
    .X(_02770_));
 sky130_fd_sc_hd__or2b_1 _10097_ (.A(_02496_),
    .B_N(_04391_),
    .X(_02771_));
 sky130_fd_sc_hd__or2b_1 _10098_ (.A(_04380_),
    .B_N(_02496_),
    .X(_02772_));
 sky130_fd_sc_hd__and2_1 _10099_ (.A(_02771_),
    .B(_02772_),
    .X(_02773_));
 sky130_fd_sc_hd__and4_1 _10100_ (.A(_02766_),
    .B(_02769_),
    .C(_02770_),
    .D(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__nand3_1 _10101_ (.A(_02757_),
    .B(_02760_),
    .C(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__and2b_1 _10102_ (.A_N(_03293_),
    .B(_05402_),
    .X(_02777_));
 sky130_fd_sc_hd__and2b_1 _10103_ (.A_N(_05402_),
    .B(_03293_),
    .X(_02778_));
 sky130_fd_sc_hd__nor2_1 _10104_ (.A(_02777_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__and2b_1 _10105_ (.A_N(_03346_),
    .B(_05467_),
    .X(_02780_));
 sky130_fd_sc_hd__or2b_1 _10106_ (.A(_05467_),
    .B_N(_03346_),
    .X(_02781_));
 sky130_fd_sc_hd__nor2b_2 _10107_ (.A(_02780_),
    .B_N(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_1 _10108_ (.A(_02779_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__and2b_1 _10109_ (.A_N(_02550_),
    .B(_04467_),
    .X(_02784_));
 sky130_fd_sc_hd__and2b_1 _10110_ (.A_N(_04467_),
    .B(_02550_),
    .X(_02785_));
 sky130_fd_sc_hd__nor2_1 _10111_ (.A(_02784_),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__or2b_1 _10112_ (.A(_04542_),
    .B_N(_02604_),
    .X(_02787_));
 sky130_fd_sc_hd__inv_2 _10113_ (.A(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__and2b_1 _10114_ (.A_N(_02604_),
    .B(_04542_),
    .X(_02789_));
 sky130_fd_sc_hd__nor2_2 _10115_ (.A(_02788_),
    .B(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_02786_),
    .B(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__and2b_1 _10117_ (.A_N(_04865_),
    .B(_02862_),
    .X(_02792_));
 sky130_fd_sc_hd__and2b_1 _10118_ (.A_N(_02862_),
    .B(_04865_),
    .X(_02793_));
 sky130_fd_sc_hd__or2_1 _10119_ (.A(_02792_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__buf_2 _10120_ (.A(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__or2b_1 _10121_ (.A(_02916_),
    .B_N(_04929_),
    .X(_02796_));
 sky130_fd_sc_hd__inv_2 _10122_ (.A(_02796_),
    .Y(_02798_));
 sky130_fd_sc_hd__and2b_1 _10123_ (.A_N(_04929_),
    .B(_02916_),
    .X(_02799_));
 sky130_fd_sc_hd__nor2_2 _10124_ (.A(_02798_),
    .B(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__inv_2 _10125_ (.A(_03152_),
    .Y(_02801_));
 sky130_fd_sc_hd__nor2_1 _10126_ (.A(_02801_),
    .B(_05273_),
    .Y(_02802_));
 sky130_fd_sc_hd__and2_1 _10127_ (.A(_02801_),
    .B(_05273_),
    .X(_02803_));
 sky130_fd_sc_hd__nor2_1 _10128_ (.A(_02802_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__clkbuf_4 _10129_ (.A(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__and2b_1 _10130_ (.A_N(_03239_),
    .B(_05338_),
    .X(_02806_));
 sky130_fd_sc_hd__or2b_1 _10131_ (.A(_05338_),
    .B_N(_03239_),
    .X(_02807_));
 sky130_fd_sc_hd__nor2b_2 _10132_ (.A(_02806_),
    .B_N(_02807_),
    .Y(_02809_));
 sky130_fd_sc_hd__and4b_1 _10133_ (.A_N(_02795_),
    .B(_02800_),
    .C(_02805_),
    .D(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__or3b_1 _10134_ (.A(_02783_),
    .B(_02791_),
    .C_N(_02810_),
    .X(_02811_));
 sky130_fd_sc_hd__and2_1 _10135_ (.A(_03842_),
    .B(_05992_),
    .X(_02812_));
 sky130_fd_sc_hd__or2_1 _10136_ (.A(_03842_),
    .B(_05992_),
    .X(_02813_));
 sky130_fd_sc_hd__and2b_1 _10137_ (.A_N(_02812_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__nand2_2 _10138_ (.A(_03615_),
    .B(_05777_),
    .Y(_02815_));
 sky130_fd_sc_hd__or2_1 _10139_ (.A(_03626_),
    .B(_05788_),
    .X(_02816_));
 sky130_fd_sc_hd__and2_2 _10140_ (.A(_02815_),
    .B(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__and2_1 _10141_ (.A(_03755_),
    .B(_05906_),
    .X(_02818_));
 sky130_fd_sc_hd__buf_2 _10142_ (.A(_02818_),
    .X(_02820_));
 sky130_fd_sc_hd__nor2_1 _10143_ (.A(_03755_),
    .B(_05917_),
    .Y(_02821_));
 sky130_fd_sc_hd__nor2_1 _10144_ (.A(_02820_),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__and2b_1 _10145_ (.A_N(_05853_),
    .B(_03680_),
    .X(_02823_));
 sky130_fd_sc_hd__and2b_1 _10146_ (.A_N(_03680_),
    .B(_05853_),
    .X(_02824_));
 sky130_fd_sc_hd__or2_1 _10147_ (.A(_02823_),
    .B(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__or4_2 _10148_ (.A(_02814_),
    .B(_02817_),
    .C(_02822_),
    .D(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__inv_2 _10149_ (.A(_03561_),
    .Y(_02827_));
 sky130_fd_sc_hd__nor2_1 _10150_ (.A(_02827_),
    .B(_05724_),
    .Y(_02828_));
 sky130_fd_sc_hd__and2_1 _10151_ (.A(_02827_),
    .B(_05724_),
    .X(_02829_));
 sky130_fd_sc_hd__or2_2 _10152_ (.A(_02828_),
    .B(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__and2_1 _10153_ (.A(_03507_),
    .B(_05671_),
    .X(_02831_));
 sky130_fd_sc_hd__nor2_1 _10154_ (.A(_03507_),
    .B(_05671_),
    .Y(_02832_));
 sky130_fd_sc_hd__nor2_2 _10155_ (.A(_02831_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__or2b_1 _10156_ (.A(_05595_),
    .B_N(_03454_),
    .X(_02834_));
 sky130_fd_sc_hd__inv_2 _10157_ (.A(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__and2b_1 _10158_ (.A_N(_03454_),
    .B(_05595_),
    .X(_02836_));
 sky130_fd_sc_hd__nor2_2 _10159_ (.A(_02835_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__and2b_1 _10160_ (.A_N(_03400_),
    .B(_05531_),
    .X(_02838_));
 sky130_fd_sc_hd__and2b_1 _10161_ (.A_N(_05531_),
    .B(_03400_),
    .X(_02839_));
 sky130_fd_sc_hd__nor2_2 _10162_ (.A(_02838_),
    .B(_02839_),
    .Y(_02841_));
 sky130_fd_sc_hd__or4bb_1 _10163_ (.A(_02830_),
    .B(_02833_),
    .C_N(_02837_),
    .D_N(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__nor2_1 _10164_ (.A(_02765_),
    .B(_04736_),
    .Y(_02843_));
 sky130_fd_sc_hd__nor2_2 _10165_ (.A(_00566_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__or2b_1 _10166_ (.A(_04800_),
    .B_N(_02808_),
    .X(_02845_));
 sky130_fd_sc_hd__and2b_1 _10167_ (.A_N(_02808_),
    .B(_04800_),
    .X(_02846_));
 sky130_fd_sc_hd__inv_2 _10168_ (.A(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__nand2_2 _10169_ (.A(_02845_),
    .B(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__or2b_1 _10170_ (.A(_05058_),
    .B_N(_03024_),
    .X(_02849_));
 sky130_fd_sc_hd__and2b_1 _10171_ (.A_N(_03024_),
    .B(_05058_),
    .X(_02850_));
 sky130_fd_sc_hd__inv_2 _10172_ (.A(_02850_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _10173_ (.A(_02849_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(_03067_),
    .B(_05134_),
    .Y(_02854_));
 sky130_fd_sc_hd__or2_1 _10175_ (.A(_03067_),
    .B(_05134_),
    .X(_02855_));
 sky130_fd_sc_hd__nand2_2 _10176_ (.A(_02854_),
    .B(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__or4b_1 _10177_ (.A(_02844_),
    .B(_02848_),
    .C(_02853_),
    .D_N(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__or2b_1 _10178_ (.A(_04607_),
    .B_N(_02669_),
    .X(_02858_));
 sky130_fd_sc_hd__or2b_1 _10179_ (.A(_02669_),
    .B_N(_04607_),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_2 _10180_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__inv_2 _10181_ (.A(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__and2b_1 _10182_ (.A_N(_02970_),
    .B(_04983_),
    .X(_02863_));
 sky130_fd_sc_hd__and2b_1 _10183_ (.A_N(_04994_),
    .B(_02970_),
    .X(_02864_));
 sky130_fd_sc_hd__nor2_2 _10184_ (.A(_02863_),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__and2b_1 _10185_ (.A_N(_05209_),
    .B(_03110_),
    .X(_02866_));
 sky130_fd_sc_hd__and2b_1 _10186_ (.A_N(_03110_),
    .B(_05209_),
    .X(_02867_));
 sky130_fd_sc_hd__nor2_2 _10187_ (.A(_02866_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__and2b_1 _10188_ (.A_N(_04671_),
    .B(_02723_),
    .X(_02869_));
 sky130_fd_sc_hd__and2b_1 _10189_ (.A_N(_02723_),
    .B(_04671_),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_2 _10190_ (.A(_02869_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__and4_1 _10191_ (.A(_02861_),
    .B(_02865_),
    .C(_02868_),
    .D(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__or4b_1 _10192_ (.A(_02826_),
    .B(_02842_),
    .C(_02857_),
    .D_N(_02872_),
    .X(_02874_));
 sky130_fd_sc_hd__inv_2 _10193_ (.A(_00789_),
    .Y(_02875_));
 sky130_fd_sc_hd__inv_2 _10194_ (.A(_02842_),
    .Y(_02876_));
 sky130_fd_sc_hd__or2b_1 _10195_ (.A(_04929_),
    .B_N(_02916_),
    .X(_02877_));
 sky130_fd_sc_hd__or2b_1 _10196_ (.A(_04671_),
    .B_N(_02723_),
    .X(_02878_));
 sky130_fd_sc_hd__or2b_1 _10197_ (.A(_04262_),
    .B_N(_02388_),
    .X(_02879_));
 sky130_fd_sc_hd__or2b_1 _10198_ (.A(_04133_),
    .B_N(_02302_),
    .X(_02880_));
 sky130_fd_sc_hd__or2b_1 _10199_ (.A(_02216_),
    .B_N(_03993_),
    .X(_02881_));
 sky130_fd_sc_hd__a21bo_1 _10200_ (.A1(_02715_),
    .A2(_02753_),
    .B1_N(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__and2b_1 _10201_ (.A_N(_02302_),
    .B(_04122_),
    .X(_02883_));
 sky130_fd_sc_hd__and2b_1 _10202_ (.A_N(_02259_),
    .B(_04057_),
    .X(_02884_));
 sky130_fd_sc_hd__a211o_1 _10203_ (.A1(_02767_),
    .A2(_02882_),
    .B1(_02883_),
    .C1(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__a311o_1 _10204_ (.A1(_02766_),
    .A2(_02880_),
    .A3(_02885_),
    .B1(_02761_),
    .C1(_02759_),
    .X(_02886_));
 sky130_fd_sc_hd__and2b_1 _10205_ (.A_N(_02442_),
    .B(_04327_),
    .X(_02887_));
 sky130_fd_sc_hd__and2b_1 _10206_ (.A_N(_02496_),
    .B(_04391_),
    .X(_02888_));
 sky130_fd_sc_hd__a311o_1 _10207_ (.A1(_02879_),
    .A2(_02886_),
    .A3(_02757_),
    .B1(_02887_),
    .C1(_02888_),
    .X(_02889_));
 sky130_fd_sc_hd__a31o_1 _10208_ (.A1(_02786_),
    .A2(_02772_),
    .A3(_02889_),
    .B1(_02784_),
    .X(_02890_));
 sky130_fd_sc_hd__a21oi_1 _10209_ (.A1(_02787_),
    .A2(_02890_),
    .B1(_02789_),
    .Y(_02891_));
 sky130_fd_sc_hd__o21ai_1 _10210_ (.A1(_02891_),
    .A2(_02860_),
    .B1(_02859_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21oi_1 _10211_ (.A1(_02878_),
    .A2(_02892_),
    .B1(_02870_),
    .Y(_02893_));
 sky130_fd_sc_hd__or2b_1 _10212_ (.A(_02765_),
    .B_N(_04736_),
    .X(_02895_));
 sky130_fd_sc_hd__o21ai_1 _10213_ (.A1(_02893_),
    .A2(_02844_),
    .B1(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__a21oi_1 _10214_ (.A1(_02845_),
    .A2(_02896_),
    .B1(_02846_),
    .Y(_02897_));
 sky130_fd_sc_hd__o21bai_1 _10215_ (.A1(_02897_),
    .A2(_02795_),
    .B1_N(_02793_),
    .Y(_02898_));
 sky130_fd_sc_hd__a21o_1 _10216_ (.A1(_02877_),
    .A2(_02898_),
    .B1(_02798_),
    .X(_02899_));
 sky130_fd_sc_hd__a21o_1 _10217_ (.A1(_02899_),
    .A2(_02865_),
    .B1(_02863_),
    .X(_02900_));
 sky130_fd_sc_hd__a21o_1 _10218_ (.A1(_02849_),
    .A2(_02900_),
    .B1(_02850_),
    .X(_02901_));
 sky130_fd_sc_hd__and2b_1 _10219_ (.A_N(_03067_),
    .B(_05134_),
    .X(_02902_));
 sky130_fd_sc_hd__a21o_1 _10220_ (.A1(_02901_),
    .A2(_02856_),
    .B1(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__o21ba_1 _10221_ (.A1(_02867_),
    .A2(_02903_),
    .B1_N(_02866_),
    .X(_02904_));
 sky130_fd_sc_hd__a21o_1 _10222_ (.A1(_02904_),
    .A2(_02804_),
    .B1(_02803_),
    .X(_02906_));
 sky130_fd_sc_hd__a21oi_1 _10223_ (.A1(_02807_),
    .A2(_02906_),
    .B1(_02806_),
    .Y(_02907_));
 sky130_fd_sc_hd__or2_2 _10224_ (.A(_02777_),
    .B(_02778_),
    .X(_02908_));
 sky130_fd_sc_hd__o21bai_1 _10225_ (.A1(_02907_),
    .A2(_02908_),
    .B1_N(_02777_),
    .Y(_02909_));
 sky130_fd_sc_hd__a21o_1 _10226_ (.A1(_02781_),
    .A2(_02909_),
    .B1(_02780_),
    .X(_02910_));
 sky130_fd_sc_hd__and2b_1 _10227_ (.A_N(_03507_),
    .B(_05671_),
    .X(_02911_));
 sky130_fd_sc_hd__o21a_1 _10228_ (.A1(_02836_),
    .A2(_02838_),
    .B1(_02834_),
    .X(_02912_));
 sky130_fd_sc_hd__or2b_1 _10229_ (.A(_05671_),
    .B_N(_03507_),
    .X(_02913_));
 sky130_fd_sc_hd__o221a_1 _10230_ (.A1(_02827_),
    .A2(_05724_),
    .B1(_02911_),
    .B2(_02912_),
    .C1(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__a211oi_4 _10231_ (.A1(_02876_),
    .A2(_02910_),
    .B1(_02914_),
    .C1(_02829_),
    .Y(_02915_));
 sky130_fd_sc_hd__inv_2 _10232_ (.A(_03755_),
    .Y(_02917_));
 sky130_fd_sc_hd__and2_1 _10233_ (.A(_02917_),
    .B(_05917_),
    .X(_02918_));
 sky130_fd_sc_hd__and2b_1 _10234_ (.A_N(_03626_),
    .B(_05788_),
    .X(_02919_));
 sky130_fd_sc_hd__or2_1 _10235_ (.A(_02917_),
    .B(_05917_),
    .X(_02920_));
 sky130_fd_sc_hd__or2b_1 _10236_ (.A(_05853_),
    .B_N(_03680_),
    .X(_02921_));
 sky130_fd_sc_hd__o211a_1 _10237_ (.A1(_02824_),
    .A2(_02919_),
    .B1(_02920_),
    .C1(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__o21bai_1 _10238_ (.A1(_02918_),
    .A2(_02922_),
    .B1_N(_02814_),
    .Y(_02923_));
 sky130_fd_sc_hd__o221ai_4 _10239_ (.A1(_03842_),
    .A2(_02875_),
    .B1(_02826_),
    .B2(_02915_),
    .C1(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__o31a_2 _10240_ (.A1(_02775_),
    .A2(_02811_),
    .A3(_02874_),
    .B1(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_4 _10241_ (.A(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__clkbuf_4 _10242_ (.A(_02926_),
    .X(_02928_));
 sky130_fd_sc_hd__a21oi_1 _10243_ (.A1(_02715_),
    .A2(_02714_),
    .B1(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__xnor2_1 _10244_ (.A(_02755_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__clkbuf_4 _10245_ (.A(_06045_),
    .X(_02931_));
 sky130_fd_sc_hd__a32o_1 _10246_ (.A1(_02216_),
    .A2(_04004_),
    .A3(_02745_),
    .B1(_02931_),
    .B2(\FuI.Integer[1] ),
    .X(_02932_));
 sky130_fd_sc_hd__a221o_1 _10247_ (.A1(\MuI.result[1] ),
    .A2(_02739_),
    .B1(_02719_),
    .B2(_04068_),
    .C1(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__and4b_1 _10248_ (.A_N(_06023_),
    .B(_02020_),
    .C(_02064_),
    .D(_02705_),
    .X(_02934_));
 sky130_fd_sc_hd__buf_2 _10249_ (.A(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_1 _10250_ (.A(_02559_),
    .B(_02753_),
    .Y(_02936_));
 sky130_fd_sc_hd__or2_1 _10251_ (.A(_02559_),
    .B(_02753_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_4 _10252_ (.A(_02730_),
    .X(_02938_));
 sky130_fd_sc_hd__a22o_1 _10253_ (.A1(_02216_),
    .A2(_03928_),
    .B1(_04004_),
    .B2(_02118_),
    .X(_02939_));
 sky130_fd_sc_hd__o211a_1 _10254_ (.A1(_02532_),
    .A2(_02559_),
    .B1(_02741_),
    .C1(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__clkbuf_4 _10255_ (.A(_02727_),
    .X(_02941_));
 sky130_fd_sc_hd__nor2_1 _10256_ (.A(_04004_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__and2b_1 _10257_ (.A_N(_02706_),
    .B(_02729_),
    .X(_02943_));
 sky130_fd_sc_hd__clkbuf_4 _10258_ (.A(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__clkbuf_4 _10259_ (.A(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__a2bb2o_1 _10260_ (.A1_N(_02708_),
    .A2_N(_02753_),
    .B1(_02945_),
    .B2(_03928_),
    .X(_02946_));
 sky130_fd_sc_hd__a2111o_1 _10261_ (.A1(\AuI.result[1] ),
    .A2(_02938_),
    .B1(_02940_),
    .C1(_02942_),
    .D1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__o21a_1 _10262_ (.A1(_02216_),
    .A2(_04004_),
    .B1(_02724_),
    .X(_02949_));
 sky130_fd_sc_hd__a311o_1 _10263_ (.A1(_02935_),
    .A2(_02936_),
    .A3(_02937_),
    .B1(_02947_),
    .C1(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__a21o_1 _10264_ (.A1(_00815_),
    .A2(_02703_),
    .B1(_00814_),
    .X(_02951_));
 sky130_fd_sc_hd__a31o_1 _10265_ (.A1(_03820_),
    .A2(_04004_),
    .A3(_00689_),
    .B1(_00687_),
    .X(_02952_));
 sky130_fd_sc_hd__nand2_1 _10266_ (.A(_00673_),
    .B(_00710_),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_4 _10267_ (.A1(_00672_),
    .A2(_00711_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_00707_),
    .B(_00708_),
    .Y(_02955_));
 sky130_fd_sc_hd__or2_1 _10269_ (.A(_00707_),
    .B(_00708_),
    .X(_02956_));
 sky130_fd_sc_hd__a21boi_4 _10270_ (.A1(_00691_),
    .A2(_02955_),
    .B1_N(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ai_2 _10271_ (.A1(_00713_),
    .A2(_00748_),
    .B1(_00746_),
    .Y(_02958_));
 sky130_fd_sc_hd__or2b_1 _10272_ (.A(_00683_),
    .B_N(_00682_),
    .X(_02960_));
 sky130_fd_sc_hd__nand3_1 _10273_ (.A(_03733_),
    .B(_04068_),
    .C(_00684_),
    .Y(_02961_));
 sky130_fd_sc_hd__a22oi_1 _10274_ (.A1(_06442_),
    .A2(_00301_),
    .B1(_00259_),
    .B2(_03550_),
    .Y(_02962_));
 sky130_fd_sc_hd__and4_1 _10275_ (.A(_06444_),
    .B(_06442_),
    .C(_00301_),
    .D(_04305_),
    .X(_02963_));
 sky130_fd_sc_hd__nor2_1 _10276_ (.A(_02962_),
    .B(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hd__clkbuf_4 _10277_ (.A(net58),
    .X(_02965_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_02965_),
    .B(_04186_),
    .Y(_02966_));
 sky130_fd_sc_hd__xnor2_1 _10279_ (.A(_02964_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__o21ba_1 _10280_ (.A1(_00677_),
    .A2(_00681_),
    .B1_N(_00679_),
    .X(_02968_));
 sky130_fd_sc_hd__xnor2_1 _10281_ (.A(_02967_),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__nand2_1 _10282_ (.A(_06429_),
    .B(_04122_),
    .Y(_02971_));
 sky130_fd_sc_hd__xor2_1 _10283_ (.A(_02969_),
    .B(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__a21oi_1 _10284_ (.A1(_02960_),
    .A2(_02961_),
    .B1(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__and3_1 _10285_ (.A(_02960_),
    .B(_02961_),
    .C(_02972_),
    .X(_02974_));
 sky130_fd_sc_hd__nor2_2 _10286_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_03798_),
    .B(_04068_),
    .Y(_02976_));
 sky130_fd_sc_hd__xnor2_4 _10288_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__a21o_1 _10289_ (.A1(_00733_),
    .A2(_00741_),
    .B1(_00740_),
    .X(_02978_));
 sky130_fd_sc_hd__o21bai_1 _10290_ (.A1(_00729_),
    .A2(_00732_),
    .B1_N(_00730_),
    .Y(_02979_));
 sky130_fd_sc_hd__buf_4 _10291_ (.A(_03432_),
    .X(_02980_));
 sky130_fd_sc_hd__a22o_1 _10292_ (.A1(_02980_),
    .A2(_00093_),
    .B1(_04520_),
    .B2(_00281_),
    .X(_02982_));
 sky130_fd_sc_hd__buf_4 _10293_ (.A(_00278_),
    .X(_02983_));
 sky130_fd_sc_hd__buf_4 _10294_ (.A(_03432_),
    .X(_02984_));
 sky130_fd_sc_hd__nand4_2 _10295_ (.A(_02983_),
    .B(_02984_),
    .C(_00093_),
    .D(_04520_),
    .Y(_02985_));
 sky130_fd_sc_hd__a22o_1 _10296_ (.A1(_00345_),
    .A2(_04380_),
    .B1(_02982_),
    .B2(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_8 _10297_ (.A(_00292_),
    .X(_02987_));
 sky130_fd_sc_hd__nand4_2 _10298_ (.A(_02987_),
    .B(_04380_),
    .C(_02982_),
    .D(_02985_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand3_2 _10299_ (.A(_02979_),
    .B(_02986_),
    .C(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__a21o_1 _10300_ (.A1(_02986_),
    .A2(_02988_),
    .B1(_02979_),
    .X(_02990_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_00695_),
    .B(_00697_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21o_1 _10302_ (.A1(_02989_),
    .A2(_02990_),
    .B1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__nand3_1 _10303_ (.A(_02991_),
    .B(_02989_),
    .C(_02990_),
    .Y(_02993_));
 sky130_fd_sc_hd__and3_1 _10304_ (.A(_02978_),
    .B(_02992_),
    .C(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__a21oi_1 _10305_ (.A1(_02992_),
    .A2(_02993_),
    .B1(_02978_),
    .Y(_02995_));
 sky130_fd_sc_hd__a211oi_1 _10306_ (.A1(_00698_),
    .A2(_00702_),
    .B1(_02994_),
    .C1(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__o211a_1 _10307_ (.A1(_02994_),
    .A2(_02995_),
    .B1(_00698_),
    .C1(_00702_),
    .X(_02997_));
 sky130_fd_sc_hd__nor2_1 _10308_ (.A(_02996_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nor2_2 _10309_ (.A(_00703_),
    .B(_00705_),
    .Y(_02999_));
 sky130_fd_sc_hd__xnor2_2 _10310_ (.A(_02998_),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__xnor2_2 _10311_ (.A(_02977_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__xor2_2 _10312_ (.A(_02958_),
    .B(_03001_),
    .X(_03003_));
 sky130_fd_sc_hd__xor2_2 _10313_ (.A(_02957_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nor2_1 _10314_ (.A(_00725_),
    .B(_00745_),
    .Y(_03005_));
 sky130_fd_sc_hd__nand3_1 _10315_ (.A(_00750_),
    .B(_00764_),
    .C(_00765_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_00716_),
    .B(_00717_),
    .Y(_03007_));
 sky130_fd_sc_hd__o21bai_1 _10317_ (.A1(_00751_),
    .A2(_00754_),
    .B1_N(_00752_),
    .Y(_03008_));
 sky130_fd_sc_hd__a22o_1 _10318_ (.A1(_02959_),
    .A2(_00421_),
    .B1(_00534_),
    .B2(_00217_),
    .X(_03009_));
 sky130_fd_sc_hd__nand4_1 _10319_ (.A(_02905_),
    .B(_02959_),
    .C(_00421_),
    .D(_00423_),
    .Y(_03010_));
 sky130_fd_sc_hd__a22o_1 _10320_ (.A1(_03013_),
    .A2(_04983_),
    .B1(_03009_),
    .B2(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__nand4_1 _10321_ (.A(_03013_),
    .B(_04983_),
    .C(_03009_),
    .D(_03010_),
    .Y(_03012_));
 sky130_fd_sc_hd__nand3_1 _10322_ (.A(_03008_),
    .B(_03011_),
    .C(_03012_),
    .Y(_03014_));
 sky130_fd_sc_hd__a21o_1 _10323_ (.A1(_03011_),
    .A2(_03012_),
    .B1(_03008_),
    .X(_03015_));
 sky130_fd_sc_hd__nand3_1 _10324_ (.A(_03007_),
    .B(_03014_),
    .C(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__a21o_1 _10325_ (.A1(_03014_),
    .A2(_03015_),
    .B1(_03007_),
    .X(_03017_));
 sky130_fd_sc_hd__a21bo_1 _10326_ (.A1(_00721_),
    .A2(_00720_),
    .B1_N(_00719_),
    .X(_03018_));
 sky130_fd_sc_hd__and3_1 _10327_ (.A(_03016_),
    .B(_03017_),
    .C(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__a21oi_1 _10328_ (.A1(_03016_),
    .A2(_03017_),
    .B1(_03018_),
    .Y(_03020_));
 sky130_fd_sc_hd__a22oi_1 _10329_ (.A1(_00727_),
    .A2(_00059_),
    .B1(_04714_),
    .B2(_00728_),
    .Y(_03021_));
 sky130_fd_sc_hd__and4_1 _10330_ (.A(_01147_),
    .B(_01146_),
    .C(_04649_),
    .D(_04714_),
    .X(_03022_));
 sky130_fd_sc_hd__nor2_1 _10331_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(_00077_),
    .B(_04596_),
    .Y(_03025_));
 sky130_fd_sc_hd__xnor2_1 _10333_ (.A(_03023_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__a22o_1 _10334_ (.A1(_01206_),
    .A2(_04843_),
    .B1(_04907_),
    .B2(_00921_),
    .X(_03027_));
 sky130_fd_sc_hd__nand4_1 _10335_ (.A(_03067_),
    .B(_01206_),
    .C(_00445_),
    .D(_00550_),
    .Y(_03028_));
 sky130_fd_sc_hd__and2_1 _10336_ (.A(_03163_),
    .B(_04789_),
    .X(_03029_));
 sky130_fd_sc_hd__a21o_1 _10337_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__nand3_1 _10338_ (.A(_03029_),
    .B(_03027_),
    .C(_03028_),
    .Y(_03031_));
 sky130_fd_sc_hd__o21bai_1 _10339_ (.A1(_00734_),
    .A2(_00736_),
    .B1_N(_00735_),
    .Y(_03032_));
 sky130_fd_sc_hd__and3_1 _10340_ (.A(_03030_),
    .B(_03031_),
    .C(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__a21o_1 _10341_ (.A1(_03030_),
    .A2(_03031_),
    .B1(_03032_),
    .X(_03034_));
 sky130_fd_sc_hd__and2b_1 _10342_ (.A_N(_03033_),
    .B(_03034_),
    .X(_03036_));
 sky130_fd_sc_hd__xnor2_1 _10343_ (.A(_03026_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__o21a_1 _10344_ (.A1(_03019_),
    .A2(_03020_),
    .B1(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__nor3_1 _10345_ (.A(_03037_),
    .B(_03019_),
    .C(_03020_),
    .Y(_03039_));
 sky130_fd_sc_hd__a211o_1 _10346_ (.A1(_03006_),
    .A2(_00768_),
    .B1(_03038_),
    .C1(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__o211ai_1 _10347_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_03006_),
    .C1(_00768_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_1 _10348_ (.A(_03040_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__xor2_2 _10349_ (.A(_03005_),
    .B(_03042_),
    .X(_03043_));
 sky130_fd_sc_hd__a21o_1 _10350_ (.A1(_00771_),
    .A2(_00779_),
    .B1(_00778_),
    .X(_03044_));
 sky130_fd_sc_hd__nand2_1 _10351_ (.A(_06610_),
    .B(_05198_),
    .Y(_03045_));
 sky130_fd_sc_hd__a22oi_4 _10352_ (.A1(_02808_),
    .A2(_05262_),
    .B1(_05327_),
    .B2(_02765_),
    .Y(_03046_));
 sky130_fd_sc_hd__buf_4 _10353_ (.A(_05305_),
    .X(_03047_));
 sky130_fd_sc_hd__and4_1 _10354_ (.A(_00877_),
    .B(_00878_),
    .C(_06561_),
    .D(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__nor2_1 _10355_ (.A(_03046_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__xnor2_1 _10356_ (.A(_03045_),
    .B(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__clkbuf_4 _10357_ (.A(_05498_),
    .X(_03051_));
 sky130_fd_sc_hd__a22o_1 _10358_ (.A1(_06682_),
    .A2(_06546_),
    .B1(_03051_),
    .B2(_00000_),
    .X(_03052_));
 sky130_fd_sc_hd__nand4_1 _10359_ (.A(_02604_),
    .B(_02669_),
    .C(_06546_),
    .D(_03051_),
    .Y(_03053_));
 sky130_fd_sc_hd__and2_1 _10360_ (.A(_06593_),
    .B(_06477_),
    .X(_03054_));
 sky130_fd_sc_hd__a21o_1 _10361_ (.A1(_03052_),
    .A2(_03053_),
    .B1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__nand3_1 _10362_ (.A(_03054_),
    .B(_03052_),
    .C(_03053_),
    .Y(_03057_));
 sky130_fd_sc_hd__o21bai_1 _10363_ (.A1(_00756_),
    .A2(_00758_),
    .B1_N(_00757_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand3_1 _10364_ (.A(_03055_),
    .B(_03057_),
    .C(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__a21o_1 _10365_ (.A1(_03055_),
    .A2(_03057_),
    .B1(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__nand3_1 _10366_ (.A(_03050_),
    .B(_03059_),
    .C(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__a21o_1 _10367_ (.A1(_03059_),
    .A2(_03060_),
    .B1(_03050_),
    .X(_03062_));
 sky130_fd_sc_hd__and3_1 _10368_ (.A(_03044_),
    .B(_03061_),
    .C(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__a21oi_1 _10369_ (.A1(_03061_),
    .A2(_03062_),
    .B1(_03044_),
    .Y(_03064_));
 sky130_fd_sc_hd__a211oi_1 _10370_ (.A1(_00762_),
    .A2(_00764_),
    .B1(_03063_),
    .C1(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__o211a_1 _10371_ (.A1(_03063_),
    .A2(_03064_),
    .B1(_00762_),
    .C1(_00764_),
    .X(_03066_));
 sky130_fd_sc_hd__nor2_1 _10372_ (.A(_03065_),
    .B(_03066_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_1 _10373_ (.A(_00774_),
    .B(_00776_),
    .Y(_03069_));
 sky130_fd_sc_hd__o21bai_1 _10374_ (.A1(_00782_),
    .A2(_00784_),
    .B1_N(_00786_),
    .Y(_03070_));
 sky130_fd_sc_hd__buf_4 _10375_ (.A(_05563_),
    .X(_03071_));
 sky130_fd_sc_hd__a22o_1 _10376_ (.A1(_02485_),
    .A2(_05638_),
    .B1(_06537_),
    .B2(_06565_),
    .X(_03072_));
 sky130_fd_sc_hd__nand4_1 _10377_ (.A(_02431_),
    .B(_02485_),
    .C(_00382_),
    .D(_00163_),
    .Y(_03073_));
 sky130_fd_sc_hd__a22o_1 _10378_ (.A1(_06560_),
    .A2(_03071_),
    .B1(_03072_),
    .B2(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__nand4_1 _10379_ (.A(_02539_),
    .B(_03071_),
    .C(_03072_),
    .D(_03073_),
    .Y(_03075_));
 sky130_fd_sc_hd__and3_1 _10380_ (.A(_03070_),
    .B(_03074_),
    .C(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__a21o_1 _10381_ (.A1(_03074_),
    .A2(_03075_),
    .B1(_03070_),
    .X(_03077_));
 sky130_fd_sc_hd__and2b_1 _10382_ (.A_N(_03076_),
    .B(_03077_),
    .X(_03079_));
 sky130_fd_sc_hd__xor2_2 _10383_ (.A(_03069_),
    .B(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__a22o_1 _10384_ (.A1(_06500_),
    .A2(_00785_),
    .B1(_00153_),
    .B2(_06501_),
    .X(_03081_));
 sky130_fd_sc_hd__buf_2 _10385_ (.A(net28),
    .X(_03082_));
 sky130_fd_sc_hd__nand4_1 _10386_ (.A(_00164_),
    .B(_00162_),
    .C(_00783_),
    .D(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__and2_1 _10387_ (.A(net108),
    .B(_05756_),
    .X(_03084_));
 sky130_fd_sc_hd__a21o_1 _10388_ (.A1(_03081_),
    .A2(_03083_),
    .B1(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__nand3_1 _10389_ (.A(_03081_),
    .B(_03083_),
    .C(_03084_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _10390_ (.A(_02216_),
    .B(_05884_),
    .Y(_03087_));
 sky130_fd_sc_hd__and3_1 _10391_ (.A(_02259_),
    .B(_05948_),
    .C(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__a21oi_1 _10392_ (.A1(_03085_),
    .A2(_03086_),
    .B1(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__and3_1 _10393_ (.A(_03085_),
    .B(_03086_),
    .C(_03088_),
    .X(_03090_));
 sky130_fd_sc_hd__or2_1 _10394_ (.A(_03089_),
    .B(_03090_),
    .X(_03091_));
 sky130_fd_sc_hd__and2b_1 _10395_ (.A_N(_00792_),
    .B(_00793_),
    .X(_03092_));
 sky130_fd_sc_hd__a21oi_2 _10396_ (.A1(_00788_),
    .A2(_00794_),
    .B1(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__xnor2_1 _10397_ (.A(_03091_),
    .B(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__xnor2_2 _10398_ (.A(_03080_),
    .B(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__or2b_1 _10399_ (.A(_00795_),
    .B_N(_00796_),
    .X(_03096_));
 sky130_fd_sc_hd__o21a_1 _10400_ (.A1(_00781_),
    .A2(_00797_),
    .B1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__xnor2_1 _10401_ (.A(_03095_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__xnor2_2 _10402_ (.A(_03068_),
    .B(_03098_),
    .Y(_03100_));
 sky130_fd_sc_hd__and2b_1 _10403_ (.A_N(_00798_),
    .B(_00799_),
    .X(_03101_));
 sky130_fd_sc_hd__a21oi_2 _10404_ (.A1(_00770_),
    .A2(_00800_),
    .B1(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__xor2_2 _10405_ (.A(_03100_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__xor2_2 _10406_ (.A(_03043_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__and2b_1 _10407_ (.A_N(_00801_),
    .B(_00802_),
    .X(_03105_));
 sky130_fd_sc_hd__a21oi_1 _10408_ (.A1(_00749_),
    .A2(_00803_),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__xnor2_2 _10409_ (.A(_03104_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__xnor2_2 _10410_ (.A(_03004_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__and2b_1 _10411_ (.A_N(_00805_),
    .B(_00804_),
    .X(_03109_));
 sky130_fd_sc_hd__a21oi_2 _10412_ (.A1(_00712_),
    .A2(_00806_),
    .B1(_03109_),
    .Y(_03111_));
 sky130_fd_sc_hd__xnor2_2 _10413_ (.A(_03108_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__xnor2_4 _10414_ (.A(_02954_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _10415_ (.A(_00807_),
    .B(_00808_),
    .Y(_03114_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_00807_),
    .B(_00808_),
    .Y(_03115_));
 sky130_fd_sc_hd__a21oi_4 _10417_ (.A1(_00669_),
    .A2(_03114_),
    .B1(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__xnor2_1 _10418_ (.A(_03113_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__xnor2_1 _10419_ (.A(_02952_),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _10420_ (.A(_00810_),
    .B(_00811_),
    .Y(_03119_));
 sky130_fd_sc_hd__a21oi_1 _10421_ (.A1(_00666_),
    .A2(_00812_),
    .B1(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(_03118_),
    .B(_03120_),
    .Y(_03122_));
 sky130_fd_sc_hd__nand2_1 _10423_ (.A(_03118_),
    .B(_03120_),
    .Y(_03123_));
 sky130_fd_sc_hd__and2b_1 _10424_ (.A_N(_03122_),
    .B(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(_02951_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__nor2_1 _10426_ (.A(_06428_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__or3_1 _10427_ (.A(_02933_),
    .B(_02950_),
    .C(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__a21o_2 _10428_ (.A1(_02752_),
    .A2(_02930_),
    .B1(_03127_),
    .X(net80));
 sky130_fd_sc_hd__xnor2_1 _10429_ (.A(_02767_),
    .B(_02882_),
    .Y(_03128_));
 sky130_fd_sc_hd__o21ai_1 _10430_ (.A1(_02770_),
    .A2(_02928_),
    .B1(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__or3_1 _10431_ (.A(_02770_),
    .B(_02928_),
    .C(_03128_),
    .X(_03130_));
 sky130_fd_sc_hd__and3_1 _10432_ (.A(_02020_),
    .B(_06023_),
    .C(_02140_),
    .X(_03132_));
 sky130_fd_sc_hd__clkbuf_4 _10433_ (.A(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__clkbuf_4 _10434_ (.A(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__a31o_1 _10435_ (.A1(_03831_),
    .A2(_04068_),
    .A3(_02975_),
    .B1(_02973_),
    .X(_03135_));
 sky130_fd_sc_hd__or2b_1 _10436_ (.A(_03001_),
    .B_N(_02958_),
    .X(_03136_));
 sky130_fd_sc_hd__o21ai_4 _10437_ (.A1(_02957_),
    .A2(_03003_),
    .B1(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__or2b_1 _10438_ (.A(_02999_),
    .B_N(_02998_),
    .X(_03138_));
 sky130_fd_sc_hd__a21boi_2 _10439_ (.A1(_02977_),
    .A2(_03000_),
    .B1_N(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__o21ai_2 _10440_ (.A1(_03005_),
    .A2(_03042_),
    .B1(_03040_),
    .Y(_03140_));
 sky130_fd_sc_hd__or2b_1 _10441_ (.A(_02968_),
    .B_N(_02967_),
    .X(_03141_));
 sky130_fd_sc_hd__nand3_1 _10442_ (.A(_03733_),
    .B(_04133_),
    .C(_02969_),
    .Y(_03142_));
 sky130_fd_sc_hd__a22oi_1 _10443_ (.A1(_03615_),
    .A2(_00259_),
    .B1(_04369_),
    .B2(_03550_),
    .Y(_03143_));
 sky130_fd_sc_hd__and4_1 _10444_ (.A(_06444_),
    .B(_06442_),
    .C(_00259_),
    .D(_04369_),
    .X(_03144_));
 sky130_fd_sc_hd__nor2_1 _10445_ (.A(_03143_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _10446_ (.A(_02965_),
    .B(_04251_),
    .Y(_03146_));
 sky130_fd_sc_hd__xnor2_1 _10447_ (.A(_03145_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__o21ba_1 _10448_ (.A1(_02962_),
    .A2(_02966_),
    .B1_N(_02963_),
    .X(_03148_));
 sky130_fd_sc_hd__xnor2_1 _10449_ (.A(_03147_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_06429_),
    .B(_04197_),
    .Y(_03150_));
 sky130_fd_sc_hd__xor2_1 _10451_ (.A(_03149_),
    .B(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__a21oi_1 _10452_ (.A1(_03141_),
    .A2(_03142_),
    .B1(_03151_),
    .Y(_03153_));
 sky130_fd_sc_hd__and3_1 _10453_ (.A(_03141_),
    .B(_03142_),
    .C(_03151_),
    .X(_03154_));
 sky130_fd_sc_hd__nor2_2 _10454_ (.A(_03153_),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_03798_),
    .B(_04133_),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_4 _10456_ (.A(_03155_),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_1 _10457_ (.A1(_03026_),
    .A2(_03034_),
    .B1(_03033_),
    .X(_03158_));
 sky130_fd_sc_hd__o21bai_1 _10458_ (.A1(_03021_),
    .A2(_03025_),
    .B1_N(_03022_),
    .Y(_03159_));
 sky130_fd_sc_hd__a22o_1 _10459_ (.A1(_02984_),
    .A2(_04520_),
    .B1(_00036_),
    .B2(_02983_),
    .X(_03160_));
 sky130_fd_sc_hd__nand4_2 _10460_ (.A(_03389_),
    .B(_02984_),
    .C(_04520_),
    .D(_00036_),
    .Y(_03161_));
 sky130_fd_sc_hd__a22o_1 _10461_ (.A1(_02987_),
    .A2(_04456_),
    .B1(_03160_),
    .B2(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__nand4_2 _10462_ (.A(_02987_),
    .B(_04456_),
    .C(_03160_),
    .D(_03161_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand3_2 _10463_ (.A(_03159_),
    .B(_03162_),
    .C(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__a21o_1 _10464_ (.A1(_03162_),
    .A2(_03164_),
    .B1(_03159_),
    .X(_03166_));
 sky130_fd_sc_hd__nand2_1 _10465_ (.A(_02985_),
    .B(_02988_),
    .Y(_03167_));
 sky130_fd_sc_hd__a21o_1 _10466_ (.A1(_03165_),
    .A2(_03166_),
    .B1(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nand3_2 _10467_ (.A(_03167_),
    .B(_03165_),
    .C(_03166_),
    .Y(_03169_));
 sky130_fd_sc_hd__and3_1 _10468_ (.A(_03158_),
    .B(_03168_),
    .C(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__a21oi_1 _10469_ (.A1(_03168_),
    .A2(_03169_),
    .B1(_03158_),
    .Y(_03171_));
 sky130_fd_sc_hd__a211oi_2 _10470_ (.A1(_02989_),
    .A2(_02993_),
    .B1(_03170_),
    .C1(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__o211a_1 _10471_ (.A1(_03170_),
    .A2(_03171_),
    .B1(_02989_),
    .C1(_02993_),
    .X(_03173_));
 sky130_fd_sc_hd__nor2_1 _10472_ (.A(_03172_),
    .B(_03173_),
    .Y(_03175_));
 sky130_fd_sc_hd__nor2_1 _10473_ (.A(_02994_),
    .B(_02996_),
    .Y(_03176_));
 sky130_fd_sc_hd__xnor2_2 _10474_ (.A(_03175_),
    .B(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__xnor2_2 _10475_ (.A(_03157_),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__xor2_2 _10476_ (.A(_03140_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__xor2_2 _10477_ (.A(_03139_),
    .B(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__nor2_1 _10478_ (.A(_03019_),
    .B(_03039_),
    .Y(_03181_));
 sky130_fd_sc_hd__o21bai_1 _10479_ (.A1(_03045_),
    .A2(_03046_),
    .B1_N(_03048_),
    .Y(_03182_));
 sky130_fd_sc_hd__a22o_1 _10480_ (.A1(_02959_),
    .A2(_00423_),
    .B1(_05198_),
    .B2(_02905_),
    .X(_03183_));
 sky130_fd_sc_hd__nand4_1 _10481_ (.A(_02905_),
    .B(_02959_),
    .C(_00423_),
    .D(_05198_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_4 _10482_ (.A(_00058_),
    .B(_00421_),
    .Y(_03186_));
 sky130_fd_sc_hd__a21bo_1 _10483_ (.A1(_03183_),
    .A2(_03184_),
    .B1_N(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__nand3b_1 _10484_ (.A_N(_03186_),
    .B(_03183_),
    .C(_03184_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand3_1 _10485_ (.A(_03182_),
    .B(_03187_),
    .C(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__a21o_1 _10486_ (.A1(_03187_),
    .A2(_03188_),
    .B1(_03182_),
    .X(_03190_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_03010_),
    .B(_03012_),
    .Y(_03191_));
 sky130_fd_sc_hd__a21o_1 _10488_ (.A1(_03189_),
    .A2(_03190_),
    .B1(_03191_),
    .X(_03192_));
 sky130_fd_sc_hd__nand3_1 _10489_ (.A(_03191_),
    .B(_03189_),
    .C(_03190_),
    .Y(_03193_));
 sky130_fd_sc_hd__a21bo_1 _10490_ (.A1(_03007_),
    .A2(_03015_),
    .B1_N(_03014_),
    .X(_03194_));
 sky130_fd_sc_hd__nand3_1 _10491_ (.A(_03192_),
    .B(_03193_),
    .C(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__a21o_1 _10492_ (.A1(_03192_),
    .A2(_03193_),
    .B1(_03194_),
    .X(_03197_));
 sky130_fd_sc_hd__a22oi_1 _10493_ (.A1(_00727_),
    .A2(_04714_),
    .B1(_06613_),
    .B2(_00728_),
    .Y(_03198_));
 sky130_fd_sc_hd__and4_1 _10494_ (.A(_01147_),
    .B(_01146_),
    .C(_04714_),
    .D(_04789_),
    .X(_03199_));
 sky130_fd_sc_hd__nor2_1 _10495_ (.A(_03198_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _10496_ (.A(_00077_),
    .B(_00059_),
    .Y(_03201_));
 sky130_fd_sc_hd__xnor2_1 _10497_ (.A(_03200_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hd__a22o_1 _10498_ (.A1(_01206_),
    .A2(_04907_),
    .B1(_04972_),
    .B2(_00921_),
    .X(_03203_));
 sky130_fd_sc_hd__nand4_1 _10499_ (.A(_00921_),
    .B(_01206_),
    .C(_04907_),
    .D(_04972_),
    .Y(_03204_));
 sky130_fd_sc_hd__and2_1 _10500_ (.A(_03163_),
    .B(_04843_),
    .X(_03205_));
 sky130_fd_sc_hd__a21o_1 _10501_ (.A1(_03203_),
    .A2(_03204_),
    .B1(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__nand3_1 _10502_ (.A(_03205_),
    .B(_03203_),
    .C(_03204_),
    .Y(_03207_));
 sky130_fd_sc_hd__a21bo_1 _10503_ (.A1(_03029_),
    .A2(_03027_),
    .B1_N(_03028_),
    .X(_03208_));
 sky130_fd_sc_hd__and3_1 _10504_ (.A(_03206_),
    .B(_03207_),
    .C(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__a21o_1 _10505_ (.A1(_03206_),
    .A2(_03207_),
    .B1(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__or2b_1 _10506_ (.A(_03209_),
    .B_N(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__xnor2_1 _10507_ (.A(_03202_),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__a21o_1 _10508_ (.A1(_03195_),
    .A2(_03197_),
    .B1(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__nand3_1 _10509_ (.A(_03212_),
    .B(_03195_),
    .C(_03197_),
    .Y(_03214_));
 sky130_fd_sc_hd__o211ai_1 _10510_ (.A1(_03063_),
    .A2(_03065_),
    .B1(_03213_),
    .C1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__a211o_1 _10511_ (.A1(_03213_),
    .A2(_03214_),
    .B1(_03063_),
    .C1(_03065_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(_03215_),
    .B(_03216_),
    .Y(_03218_));
 sky130_fd_sc_hd__xor2_1 _10513_ (.A(_03181_),
    .B(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__nand2_1 _10514_ (.A(_03059_),
    .B(_03061_),
    .Y(_03220_));
 sky130_fd_sc_hd__a21o_1 _10515_ (.A1(_03069_),
    .A2(_03077_),
    .B1(_03076_),
    .X(_03221_));
 sky130_fd_sc_hd__nand2_1 _10516_ (.A(_02840_),
    .B(_06561_),
    .Y(_03222_));
 sky130_fd_sc_hd__a22oi_1 _10517_ (.A1(_02808_),
    .A2(_03047_),
    .B1(_06477_),
    .B2(_02765_),
    .Y(_03223_));
 sky130_fd_sc_hd__and4_1 _10518_ (.A(_06606_),
    .B(_06601_),
    .C(_05316_),
    .D(_05380_),
    .X(_03224_));
 sky130_fd_sc_hd__nor2_1 _10519_ (.A(_03223_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__xnor2_1 _10520_ (.A(_03222_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__a22o_1 _10521_ (.A1(_06682_),
    .A2(_05509_),
    .B1(_05574_),
    .B2(_00000_),
    .X(_03227_));
 sky130_fd_sc_hd__nand4_1 _10522_ (.A(_00000_),
    .B(_02669_),
    .C(_03051_),
    .D(_03071_),
    .Y(_03229_));
 sky130_fd_sc_hd__and2_1 _10523_ (.A(_06593_),
    .B(_05445_),
    .X(_03230_));
 sky130_fd_sc_hd__a21o_1 _10524_ (.A1(_03227_),
    .A2(_03229_),
    .B1(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__nand3_1 _10525_ (.A(_03230_),
    .B(_03227_),
    .C(_03229_),
    .Y(_03232_));
 sky130_fd_sc_hd__a21bo_1 _10526_ (.A1(_03054_),
    .A2(_03052_),
    .B1_N(_03053_),
    .X(_03233_));
 sky130_fd_sc_hd__nand3_1 _10527_ (.A(_03231_),
    .B(_03232_),
    .C(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__a21o_1 _10528_ (.A1(_03231_),
    .A2(_03232_),
    .B1(_03233_),
    .X(_03235_));
 sky130_fd_sc_hd__nand3_1 _10529_ (.A(_03226_),
    .B(_03234_),
    .C(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__a21o_1 _10530_ (.A1(_03234_),
    .A2(_03235_),
    .B1(_03226_),
    .X(_03237_));
 sky130_fd_sc_hd__nand3_1 _10531_ (.A(_03221_),
    .B(_03236_),
    .C(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__a21o_1 _10532_ (.A1(_03236_),
    .A2(_03237_),
    .B1(_03221_),
    .X(_03240_));
 sky130_fd_sc_hd__and3_1 _10533_ (.A(_03220_),
    .B(_03238_),
    .C(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__a21oi_1 _10534_ (.A1(_03238_),
    .A2(_03240_),
    .B1(_03220_),
    .Y(_03242_));
 sky130_fd_sc_hd__nor2_1 _10535_ (.A(_03241_),
    .B(_03242_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand2_1 _10536_ (.A(_03073_),
    .B(_03075_),
    .Y(_03244_));
 sky130_fd_sc_hd__a21bo_1 _10537_ (.A1(_03081_),
    .A2(_03084_),
    .B1_N(_03083_),
    .X(_03245_));
 sky130_fd_sc_hd__a22o_1 _10538_ (.A1(_02229_),
    .A2(_06537_),
    .B1(_00385_),
    .B2(_02431_),
    .X(_03246_));
 sky130_fd_sc_hd__clkbuf_4 _10539_ (.A(net25),
    .X(_03247_));
 sky130_fd_sc_hd__nand4_1 _10540_ (.A(_02431_),
    .B(_02229_),
    .C(_00163_),
    .D(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__a22o_1 _10541_ (.A1(_06560_),
    .A2(_05649_),
    .B1(_03246_),
    .B2(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__nand4_1 _10542_ (.A(_02539_),
    .B(_05649_),
    .C(_03246_),
    .D(_03248_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand3_1 _10543_ (.A(_03245_),
    .B(_03249_),
    .C(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__a21o_1 _10544_ (.A1(_03249_),
    .A2(_03251_),
    .B1(_03245_),
    .X(_03253_));
 sky130_fd_sc_hd__nand3_1 _10545_ (.A(_03244_),
    .B(_03252_),
    .C(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__a21o_1 _10546_ (.A1(_03252_),
    .A2(_03253_),
    .B1(_03244_),
    .X(_03255_));
 sky130_fd_sc_hd__and2_1 _10547_ (.A(_03254_),
    .B(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__clkbuf_4 _10548_ (.A(_00785_),
    .X(_03257_));
 sky130_fd_sc_hd__nand2_1 _10549_ (.A(_06545_),
    .B(_03257_),
    .Y(_03258_));
 sky130_fd_sc_hd__and3_1 _10550_ (.A(_00164_),
    .B(_06500_),
    .C(_03082_),
    .X(_03259_));
 sky130_fd_sc_hd__a22o_1 _10551_ (.A1(_00162_),
    .A2(_03082_),
    .B1(_00789_),
    .B2(_00164_),
    .X(_03260_));
 sky130_fd_sc_hd__a21bo_1 _10552_ (.A1(_05948_),
    .A2(_03259_),
    .B1_N(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__xor2_1 _10553_ (.A(_03258_),
    .B(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__o21a_1 _10554_ (.A1(_00791_),
    .A2(_03090_),
    .B1(_03262_),
    .X(_03263_));
 sky130_fd_sc_hd__or3_1 _10555_ (.A(_00791_),
    .B(_03090_),
    .C(_03262_),
    .X(_03264_));
 sky130_fd_sc_hd__and2b_1 _10556_ (.A_N(_03263_),
    .B(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__xnor2_2 _10557_ (.A(_03256_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(_03091_),
    .B(_03093_),
    .Y(_03267_));
 sky130_fd_sc_hd__nor2_1 _10559_ (.A(_03091_),
    .B(_03093_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21oi_2 _10560_ (.A1(_03080_),
    .A2(_03267_),
    .B1(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__xor2_2 _10561_ (.A(_03266_),
    .B(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__xnor2_2 _10562_ (.A(_03243_),
    .B(_03270_),
    .Y(_03272_));
 sky130_fd_sc_hd__and2b_1 _10563_ (.A_N(_03097_),
    .B(_03095_),
    .X(_03273_));
 sky130_fd_sc_hd__a21oi_1 _10564_ (.A1(_03068_),
    .A2(_03098_),
    .B1(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__xor2_1 _10565_ (.A(_03272_),
    .B(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__xor2_1 _10566_ (.A(_03219_),
    .B(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__nor2_1 _10567_ (.A(_03100_),
    .B(_03102_),
    .Y(_03277_));
 sky130_fd_sc_hd__a21oi_1 _10568_ (.A1(_03043_),
    .A2(_03103_),
    .B1(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__xnor2_1 _10569_ (.A(_03276_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__xnor2_2 _10570_ (.A(_03180_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__and2b_1 _10571_ (.A_N(_03106_),
    .B(_03104_),
    .X(_03281_));
 sky130_fd_sc_hd__a21oi_2 _10572_ (.A1(_03004_),
    .A2(_03107_),
    .B1(_03281_),
    .Y(_03283_));
 sky130_fd_sc_hd__xnor2_2 _10573_ (.A(_03280_),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor2_4 _10574_ (.A(_03137_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _10575_ (.A(_03108_),
    .B(_03111_),
    .Y(_03286_));
 sky130_fd_sc_hd__nor2_1 _10576_ (.A(_03108_),
    .B(_03111_),
    .Y(_03287_));
 sky130_fd_sc_hd__a21oi_2 _10577_ (.A1(_02954_),
    .A2(_03286_),
    .B1(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__xnor2_4 _10578_ (.A(_03285_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__xnor2_2 _10579_ (.A(_03135_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__and2b_1 _10580_ (.A_N(_03116_),
    .B(_03113_),
    .X(_03291_));
 sky130_fd_sc_hd__a21oi_1 _10581_ (.A1(_02952_),
    .A2(_03117_),
    .B1(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__xnor2_1 _10582_ (.A(_03290_),
    .B(_03292_),
    .Y(_03294_));
 sky130_fd_sc_hd__and2b_1 _10583_ (.A_N(_00816_),
    .B(_03124_),
    .X(_03295_));
 sky130_fd_sc_hd__o21a_1 _10584_ (.A1(_00814_),
    .A2(_03122_),
    .B1(_03123_),
    .X(_03296_));
 sky130_fd_sc_hd__a21oi_1 _10585_ (.A1(_02703_),
    .A2(_03295_),
    .B1(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand2_1 _10586_ (.A(_03294_),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__or2_1 _10587_ (.A(_03294_),
    .B(_03297_),
    .X(_03299_));
 sky130_fd_sc_hd__o21ai_1 _10588_ (.A1(_02558_),
    .A2(_02560_),
    .B1(_02741_),
    .Y(_03300_));
 sky130_fd_sc_hd__nor2_1 _10589_ (.A(_02562_),
    .B(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hd__o21a_1 _10590_ (.A1(_02559_),
    .A2(_02753_),
    .B1(_02532_),
    .X(_03302_));
 sky130_fd_sc_hd__a21oi_1 _10591_ (.A1(_02767_),
    .A2(_03302_),
    .B1(_02711_),
    .Y(_03303_));
 sky130_fd_sc_hd__o21a_1 _10592_ (.A1(_02767_),
    .A2(_03302_),
    .B1(_03303_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_4 _10593_ (.A(_02720_),
    .X(_03306_));
 sky130_fd_sc_hd__o22ai_1 _10594_ (.A1(_04068_),
    .A2(_02727_),
    .B1(_02767_),
    .B2(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a221o_1 _10595_ (.A1(\MuI.result[2] ),
    .A2(_02737_),
    .B1(_02945_),
    .B2(_04004_),
    .C1(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__a32o_1 _10596_ (.A1(_02259_),
    .A2(_04068_),
    .A3(_02743_),
    .B1(_06045_),
    .B2(\FuI.Integer[2] ),
    .X(_03309_));
 sky130_fd_sc_hd__a221o_1 _10597_ (.A1(_04133_),
    .A2(_02718_),
    .B1(_02721_),
    .B2(_02259_),
    .C1(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__a211o_1 _10598_ (.A1(\AuI.result[2] ),
    .A2(_02732_),
    .B1(_03308_),
    .C1(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__or3_1 _10599_ (.A(_03301_),
    .B(_03305_),
    .C(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__a31o_1 _10600_ (.A1(_03134_),
    .A2(_03298_),
    .A3(_03299_),
    .B1(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__a31o_2 _10601_ (.A1(_02752_),
    .A2(_03129_),
    .A3(_03130_),
    .B1(_03313_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 _10602_ (.A(_02741_),
    .X(_03314_));
 sky130_fd_sc_hd__buf_4 _10603_ (.A(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__or2_1 _10604_ (.A(_02556_),
    .B(_02562_),
    .X(_03316_));
 sky130_fd_sc_hd__and2b_1 _10605_ (.A_N(_04122_),
    .B(_02302_),
    .X(_03317_));
 sky130_fd_sc_hd__or2_1 _10606_ (.A(_03317_),
    .B(_02883_),
    .X(_03318_));
 sky130_fd_sc_hd__inv_2 _10607_ (.A(_02884_),
    .Y(_03319_));
 sky130_fd_sc_hd__and2b_1 _10608_ (.A_N(_03993_),
    .B(_02216_),
    .X(_03320_));
 sky130_fd_sc_hd__a21o_1 _10609_ (.A1(_02714_),
    .A2(_02881_),
    .B1(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__and2b_1 _10610_ (.A_N(_04068_),
    .B(_02259_),
    .X(_03322_));
 sky130_fd_sc_hd__a21o_1 _10611_ (.A1(_03319_),
    .A2(_03321_),
    .B1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__a21o_1 _10612_ (.A1(_02767_),
    .A2(_02882_),
    .B1(_02884_),
    .X(_03325_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(_03323_),
    .A1(_03325_),
    .S(_02926_),
    .X(_03326_));
 sky130_fd_sc_hd__xnor2_1 _10614_ (.A(_03318_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__nor2_1 _10615_ (.A(_03290_),
    .B(_03292_),
    .Y(_03328_));
 sky130_fd_sc_hd__and2b_1 _10616_ (.A_N(_03328_),
    .B(_03299_),
    .X(_03329_));
 sky130_fd_sc_hd__and2b_2 _10617_ (.A_N(_03288_),
    .B(_03285_),
    .X(_03330_));
 sky130_fd_sc_hd__a21oi_2 _10618_ (.A1(_03135_),
    .A2(_03289_),
    .B1(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__a31o_1 _10619_ (.A1(_03820_),
    .A2(_04133_),
    .A3(_03155_),
    .B1(_03153_),
    .X(_03332_));
 sky130_fd_sc_hd__or2b_1 _10620_ (.A(_03178_),
    .B_N(_03140_),
    .X(_03333_));
 sky130_fd_sc_hd__o21ai_2 _10621_ (.A1(_03139_),
    .A2(_03179_),
    .B1(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__or2b_1 _10622_ (.A(_03176_),
    .B_N(_03175_),
    .X(_03336_));
 sky130_fd_sc_hd__a21boi_2 _10623_ (.A1(_03157_),
    .A2(_03177_),
    .B1_N(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__o21ai_2 _10624_ (.A1(_03181_),
    .A2(_03218_),
    .B1(_03215_),
    .Y(_03338_));
 sky130_fd_sc_hd__or2b_1 _10625_ (.A(_03148_),
    .B_N(_03147_),
    .X(_03339_));
 sky130_fd_sc_hd__nand3_1 _10626_ (.A(_03744_),
    .B(_04197_),
    .C(_03149_),
    .Y(_03340_));
 sky130_fd_sc_hd__a22oi_1 _10627_ (.A1(_03615_),
    .A2(_04369_),
    .B1(_04456_),
    .B2(_03550_),
    .Y(_03341_));
 sky130_fd_sc_hd__and4_1 _10628_ (.A(_06444_),
    .B(_00676_),
    .C(_00090_),
    .D(_00093_),
    .X(_03342_));
 sky130_fd_sc_hd__nor2_1 _10629_ (.A(_03341_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _10630_ (.A(_02965_),
    .B(_04316_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_1 _10631_ (.A(_03343_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21ba_1 _10632_ (.A1(_03143_),
    .A2(_03146_),
    .B1_N(_03144_),
    .X(_03347_));
 sky130_fd_sc_hd__xnor2_1 _10633_ (.A(_03345_),
    .B(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_1 _10634_ (.A(_06429_),
    .B(_04251_),
    .Y(_03349_));
 sky130_fd_sc_hd__xor2_1 _10635_ (.A(_03348_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__a21oi_1 _10636_ (.A1(_03339_),
    .A2(_03340_),
    .B1(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__and3_1 _10637_ (.A(_03339_),
    .B(_03340_),
    .C(_03350_),
    .X(_03352_));
 sky130_fd_sc_hd__nor2_2 _10638_ (.A(_03351_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_1 _10639_ (.A(_03798_),
    .B(_04197_),
    .Y(_03354_));
 sky130_fd_sc_hd__xnor2_4 _10640_ (.A(_03353_),
    .B(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hd__a21o_1 _10641_ (.A1(_03202_),
    .A2(_03210_),
    .B1(_03209_),
    .X(_03356_));
 sky130_fd_sc_hd__o21bai_1 _10642_ (.A1(_03198_),
    .A2(_03201_),
    .B1_N(_03199_),
    .Y(_03358_));
 sky130_fd_sc_hd__a22o_1 _10643_ (.A1(_02980_),
    .A2(_00036_),
    .B1(_04649_),
    .B2(_02983_),
    .X(_03359_));
 sky130_fd_sc_hd__nand4_1 _10644_ (.A(_03389_),
    .B(_02984_),
    .C(_00036_),
    .D(_00059_),
    .Y(_03360_));
 sky130_fd_sc_hd__a22o_1 _10645_ (.A1(_00345_),
    .A2(_04531_),
    .B1(_03359_),
    .B2(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__nand4_1 _10646_ (.A(_02987_),
    .B(_04531_),
    .C(_03359_),
    .D(_03360_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand3_2 _10647_ (.A(_03358_),
    .B(_03361_),
    .C(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__a21o_1 _10648_ (.A1(_03361_),
    .A2(_03362_),
    .B1(_03358_),
    .X(_03364_));
 sky130_fd_sc_hd__nand2_1 _10649_ (.A(_03161_),
    .B(_03164_),
    .Y(_03365_));
 sky130_fd_sc_hd__a21o_1 _10650_ (.A1(_03363_),
    .A2(_03364_),
    .B1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__nand3_1 _10651_ (.A(_03365_),
    .B(_03363_),
    .C(_03364_),
    .Y(_03367_));
 sky130_fd_sc_hd__and3_1 _10652_ (.A(_03356_),
    .B(_03366_),
    .C(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__a21oi_1 _10653_ (.A1(_03366_),
    .A2(_03367_),
    .B1(_03356_),
    .Y(_03369_));
 sky130_fd_sc_hd__a211o_1 _10654_ (.A1(_03165_),
    .A2(_03169_),
    .B1(_03368_),
    .C1(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__o211ai_1 _10655_ (.A1(_03368_),
    .A2(_03369_),
    .B1(_03165_),
    .C1(_03169_),
    .Y(_03371_));
 sky130_fd_sc_hd__o211ai_1 _10656_ (.A1(_03170_),
    .A2(_03172_),
    .B1(_03370_),
    .C1(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__a211o_1 _10657_ (.A1(_03370_),
    .A2(_03371_),
    .B1(_03170_),
    .C1(_03172_),
    .X(_03373_));
 sky130_fd_sc_hd__nand2_1 _10658_ (.A(_03372_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__xor2_2 _10659_ (.A(_03355_),
    .B(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__xor2_2 _10660_ (.A(_03338_),
    .B(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__xor2_1 _10661_ (.A(_03337_),
    .B(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__nand2_1 _10662_ (.A(_03195_),
    .B(_03214_),
    .Y(_03379_));
 sky130_fd_sc_hd__a31o_1 _10663_ (.A1(_03221_),
    .A2(_03236_),
    .A3(_03237_),
    .B1(_03241_),
    .X(_03380_));
 sky130_fd_sc_hd__o21bai_1 _10664_ (.A1(_03222_),
    .A2(_03223_),
    .B1_N(_03224_),
    .Y(_03381_));
 sky130_fd_sc_hd__a22o_1 _10665_ (.A1(_00062_),
    .A2(_06525_),
    .B1(_06568_),
    .B2(_00063_),
    .X(_03382_));
 sky130_fd_sc_hd__nand4_1 _10666_ (.A(_00217_),
    .B(_00216_),
    .C(_00002_),
    .D(_06568_),
    .Y(_03383_));
 sky130_fd_sc_hd__a22o_1 _10667_ (.A1(_00444_),
    .A2(_05123_),
    .B1(_03382_),
    .B2(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__nand4_1 _10668_ (.A(_00221_),
    .B(_05123_),
    .C(_03382_),
    .D(_03383_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand3_1 _10669_ (.A(_03381_),
    .B(_03384_),
    .C(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__a21o_1 _10670_ (.A1(_03384_),
    .A2(_03385_),
    .B1(_03381_),
    .X(_03387_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_03184_),
    .B(_03188_),
    .Y(_03388_));
 sky130_fd_sc_hd__a21o_1 _10672_ (.A1(_03386_),
    .A2(_03387_),
    .B1(_03388_),
    .X(_03390_));
 sky130_fd_sc_hd__nand3_1 _10673_ (.A(_03388_),
    .B(_03386_),
    .C(_03387_),
    .Y(_03391_));
 sky130_fd_sc_hd__a21bo_1 _10674_ (.A1(_03191_),
    .A2(_03190_),
    .B1_N(_03189_),
    .X(_03392_));
 sky130_fd_sc_hd__nand3_2 _10675_ (.A(_03390_),
    .B(_03391_),
    .C(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__a21o_1 _10676_ (.A1(_03390_),
    .A2(_03391_),
    .B1(_03392_),
    .X(_03394_));
 sky130_fd_sc_hd__a22oi_1 _10677_ (.A1(_00727_),
    .A2(_04789_),
    .B1(_00445_),
    .B2(_00728_),
    .Y(_03395_));
 sky130_fd_sc_hd__and4_1 _10678_ (.A(_03228_),
    .B(_03282_),
    .C(_06612_),
    .D(_04843_),
    .X(_03396_));
 sky130_fd_sc_hd__nor2_1 _10679_ (.A(_03395_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _10680_ (.A(_03324_),
    .B(_04714_),
    .Y(_03398_));
 sky130_fd_sc_hd__xnor2_1 _10681_ (.A(_03397_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__a22o_1 _10682_ (.A1(_03099_),
    .A2(_04961_),
    .B1(_06584_),
    .B2(_03056_),
    .X(_03401_));
 sky130_fd_sc_hd__nand4_1 _10683_ (.A(_00133_),
    .B(_00132_),
    .C(_06591_),
    .D(_06584_),
    .Y(_03402_));
 sky130_fd_sc_hd__and2_1 _10684_ (.A(_03152_),
    .B(_06605_),
    .X(_03403_));
 sky130_fd_sc_hd__a21o_1 _10685_ (.A1(_03401_),
    .A2(_03402_),
    .B1(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__nand3_1 _10686_ (.A(_03403_),
    .B(_03401_),
    .C(_03402_),
    .Y(_03405_));
 sky130_fd_sc_hd__a21bo_1 _10687_ (.A1(_03205_),
    .A2(_03203_),
    .B1_N(_03204_),
    .X(_03406_));
 sky130_fd_sc_hd__and3_1 _10688_ (.A(_03404_),
    .B(_03405_),
    .C(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__a21o_1 _10689_ (.A1(_03404_),
    .A2(_03405_),
    .B1(_03406_),
    .X(_03408_));
 sky130_fd_sc_hd__and2b_1 _10690_ (.A_N(_03407_),
    .B(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__xor2_1 _10691_ (.A(_03399_),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__a21o_1 _10692_ (.A1(_03393_),
    .A2(_03394_),
    .B1(_03410_),
    .X(_03412_));
 sky130_fd_sc_hd__nand3_2 _10693_ (.A(_03410_),
    .B(_03393_),
    .C(_03394_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _10694_ (.A(_03412_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _10695_ (.A(_03380_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__xor2_1 _10696_ (.A(_03379_),
    .B(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_03234_),
    .B(_03236_),
    .Y(_03417_));
 sky130_fd_sc_hd__a21bo_1 _10698_ (.A1(_03244_),
    .A2(_03253_),
    .B1_N(_03252_),
    .X(_03418_));
 sky130_fd_sc_hd__nand2_1 _10699_ (.A(net121),
    .B(_03047_),
    .Y(_03419_));
 sky130_fd_sc_hd__a22oi_1 _10700_ (.A1(_06630_),
    .A2(_05380_),
    .B1(_06546_),
    .B2(_00012_),
    .Y(_03420_));
 sky130_fd_sc_hd__and4_1 _10701_ (.A(_06598_),
    .B(_06599_),
    .C(_06476_),
    .D(_06489_),
    .X(_03421_));
 sky130_fd_sc_hd__nor2_1 _10702_ (.A(_03420_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__xnor2_1 _10703_ (.A(_03419_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__clkbuf_4 _10704_ (.A(_06461_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_4 _10705_ (.A(_05627_),
    .X(_03425_));
 sky130_fd_sc_hd__a22o_1 _10706_ (.A1(_06682_),
    .A2(_03424_),
    .B1(_03425_),
    .B2(_00000_),
    .X(_03426_));
 sky130_fd_sc_hd__nand4_1 _10707_ (.A(_00000_),
    .B(_06682_),
    .C(_05574_),
    .D(_03425_),
    .Y(_03427_));
 sky130_fd_sc_hd__and2_1 _10708_ (.A(_06680_),
    .B(_00398_),
    .X(_03428_));
 sky130_fd_sc_hd__a21o_1 _10709_ (.A1(_03426_),
    .A2(_03427_),
    .B1(_03428_),
    .X(_03429_));
 sky130_fd_sc_hd__nand3_1 _10710_ (.A(_03428_),
    .B(_03426_),
    .C(_03427_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21bo_1 _10711_ (.A1(_03230_),
    .A2(_03227_),
    .B1_N(_03229_),
    .X(_03431_));
 sky130_fd_sc_hd__nand3_1 _10712_ (.A(_03429_),
    .B(_03430_),
    .C(_03431_),
    .Y(_03433_));
 sky130_fd_sc_hd__a21o_1 _10713_ (.A1(_03429_),
    .A2(_03430_),
    .B1(_03431_),
    .X(_03434_));
 sky130_fd_sc_hd__nand3_1 _10714_ (.A(_03423_),
    .B(_03433_),
    .C(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__a21o_1 _10715_ (.A1(_03433_),
    .A2(_03434_),
    .B1(_03423_),
    .X(_03436_));
 sky130_fd_sc_hd__nand3_2 _10716_ (.A(_03418_),
    .B(_03435_),
    .C(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__a21o_1 _10717_ (.A1(_03435_),
    .A2(_03436_),
    .B1(_03418_),
    .X(_03438_));
 sky130_fd_sc_hd__nand3_2 _10718_ (.A(_03417_),
    .B(_03437_),
    .C(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__a21o_1 _10719_ (.A1(_03437_),
    .A2(_03438_),
    .B1(_03417_),
    .X(_03440_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_03439_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__a22oi_1 _10721_ (.A1(_02388_),
    .A2(_05895_),
    .B1(_05970_),
    .B2(_02345_),
    .Y(_03442_));
 sky130_fd_sc_hd__clkbuf_4 _10722_ (.A(_00153_),
    .X(_03444_));
 sky130_fd_sc_hd__and4_1 _10723_ (.A(_02345_),
    .B(_02377_),
    .C(_03444_),
    .D(_05948_),
    .X(_03445_));
 sky130_fd_sc_hd__nor2_1 _10724_ (.A(_03442_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _10725_ (.A(_03248_),
    .B(_03251_),
    .Y(_03447_));
 sky130_fd_sc_hd__a32o_1 _10726_ (.A1(_06545_),
    .A2(_03257_),
    .A3(_03260_),
    .B1(_03259_),
    .B2(_05959_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_8 _10727_ (.A(_06537_),
    .X(_03449_));
 sky130_fd_sc_hd__nand2_1 _10728_ (.A(_06560_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__nand4_1 _10729_ (.A(_02431_),
    .B(_02229_),
    .C(_03247_),
    .D(_05820_),
    .Y(_03451_));
 sky130_fd_sc_hd__a22o_1 _10730_ (.A1(_02229_),
    .A2(_00385_),
    .B1(_05820_),
    .B2(_02431_),
    .X(_03452_));
 sky130_fd_sc_hd__nand3b_1 _10731_ (.A_N(_03450_),
    .B(_03451_),
    .C(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a21bo_1 _10732_ (.A1(_03452_),
    .A2(_03451_),
    .B1_N(_03450_),
    .X(_03455_));
 sky130_fd_sc_hd__nand3_1 _10733_ (.A(_03448_),
    .B(_03453_),
    .C(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hd__a21o_1 _10734_ (.A1(_03453_),
    .A2(_03455_),
    .B1(_03448_),
    .X(_03457_));
 sky130_fd_sc_hd__nand3_1 _10735_ (.A(_03447_),
    .B(_03456_),
    .C(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21o_1 _10736_ (.A1(_03456_),
    .A2(_03457_),
    .B1(_03447_),
    .X(_03459_));
 sky130_fd_sc_hd__nand3_2 _10737_ (.A(_03446_),
    .B(_03458_),
    .C(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21o_1 _10738_ (.A1(_03458_),
    .A2(_03459_),
    .B1(_03446_),
    .X(_03461_));
 sky130_fd_sc_hd__a31o_1 _10739_ (.A1(_03254_),
    .A2(_03255_),
    .A3(_03264_),
    .B1(_03263_),
    .X(_03462_));
 sky130_fd_sc_hd__nand3_1 _10740_ (.A(_03460_),
    .B(_03461_),
    .C(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__a21o_1 _10741_ (.A1(_03460_),
    .A2(_03461_),
    .B1(_03462_),
    .X(_03464_));
 sky130_fd_sc_hd__nand2_1 _10742_ (.A(_03463_),
    .B(_03464_),
    .Y(_03466_));
 sky130_fd_sc_hd__xor2_2 _10743_ (.A(_03441_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__nor2_1 _10744_ (.A(_03266_),
    .B(_03269_),
    .Y(_03468_));
 sky130_fd_sc_hd__a21oi_1 _10745_ (.A1(_03243_),
    .A2(_03270_),
    .B1(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__xnor2_1 _10746_ (.A(_03467_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__xor2_1 _10747_ (.A(_03416_),
    .B(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__nor2_1 _10748_ (.A(_03272_),
    .B(_03274_),
    .Y(_03472_));
 sky130_fd_sc_hd__a21oi_1 _10749_ (.A1(_03219_),
    .A2(_03275_),
    .B1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__xnor2_1 _10750_ (.A(_03471_),
    .B(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__xnor2_1 _10751_ (.A(_03377_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__and2b_1 _10752_ (.A_N(_03278_),
    .B(_03276_),
    .X(_03476_));
 sky130_fd_sc_hd__a21oi_1 _10753_ (.A1(_03180_),
    .A2(_03279_),
    .B1(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__xnor2_2 _10754_ (.A(_03475_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__xnor2_2 _10755_ (.A(_03334_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(_03280_),
    .B(_03283_),
    .Y(_03480_));
 sky130_fd_sc_hd__nor2_1 _10757_ (.A(_03280_),
    .B(_03283_),
    .Y(_03481_));
 sky130_fd_sc_hd__a21oi_4 _10758_ (.A1(_03137_),
    .A2(_03480_),
    .B1(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__xnor2_4 _10759_ (.A(_03479_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__xnor2_1 _10760_ (.A(_03332_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__xnor2_1 _10761_ (.A(_03331_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(_03329_),
    .B(_03485_),
    .Y(_03487_));
 sky130_fd_sc_hd__o21a_1 _10763_ (.A1(_03329_),
    .A2(_03485_),
    .B1(_03133_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_4 _10764_ (.A(_02935_),
    .X(_03489_));
 sky130_fd_sc_hd__o21ai_1 _10765_ (.A1(_02767_),
    .A2(_03302_),
    .B1(_02498_),
    .Y(_03490_));
 sky130_fd_sc_hd__xnor2_1 _10766_ (.A(_02768_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__o21a_1 _10767_ (.A1(_02302_),
    .A2(_04133_),
    .B1(_02721_),
    .X(_03492_));
 sky130_fd_sc_hd__a221o_1 _10768_ (.A1(_02351_),
    .A2(_02745_),
    .B1(_02945_),
    .B2(_04068_),
    .C1(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__nor2_1 _10769_ (.A(_02129_),
    .B(_03306_),
    .Y(_03494_));
 sky130_fd_sc_hd__nor2_1 _10770_ (.A(_04133_),
    .B(_02726_),
    .Y(_03495_));
 sky130_fd_sc_hd__a221o_1 _10771_ (.A1(_04197_),
    .A2(_02717_),
    .B1(_02730_),
    .B2(\AuI.result[3] ),
    .C1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__a22o_1 _10772_ (.A1(\MuI.result[3] ),
    .A2(_02737_),
    .B1(_06045_),
    .B2(\FuI.Integer[3] ),
    .X(_03498_));
 sky130_fd_sc_hd__a211o_1 _10773_ (.A1(_03494_),
    .A2(_03318_),
    .B1(_03496_),
    .C1(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__or2_1 _10774_ (.A(_03493_),
    .B(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__a21o_1 _10775_ (.A1(_03489_),
    .A2(_03491_),
    .B1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__a221o_1 _10776_ (.A1(_02750_),
    .A2(_03327_),
    .B1(_03487_),
    .B2(_03488_),
    .C1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__a31o_4 _10777_ (.A1(_02563_),
    .A2(_03315_),
    .A3(_03316_),
    .B1(_03502_),
    .X(net94));
 sky130_fd_sc_hd__nand2_1 _10778_ (.A(_02880_),
    .B(_02885_),
    .Y(_03503_));
 sky130_fd_sc_hd__xnor2_1 _10779_ (.A(_02764_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__a21o_1 _10780_ (.A1(_02769_),
    .A2(_02770_),
    .B1(_02928_),
    .X(_03505_));
 sky130_fd_sc_hd__or2_1 _10781_ (.A(_03504_),
    .B(_03505_),
    .X(_03506_));
 sky130_fd_sc_hd__nand2_1 _10782_ (.A(_03504_),
    .B(_03505_),
    .Y(_03508_));
 sky130_fd_sc_hd__or2b_4 _10783_ (.A(_03482_),
    .B_N(_03479_),
    .X(_03509_));
 sky130_fd_sc_hd__nand2_1 _10784_ (.A(_03332_),
    .B(_03483_),
    .Y(_03510_));
 sky130_fd_sc_hd__a31o_1 _10785_ (.A1(_03831_),
    .A2(_04197_),
    .A3(_03353_),
    .B1(_03351_),
    .X(_03511_));
 sky130_fd_sc_hd__or2b_1 _10786_ (.A(_03375_),
    .B_N(_03338_),
    .X(_03512_));
 sky130_fd_sc_hd__o21ai_4 _10787_ (.A1(_03337_),
    .A2(_03376_),
    .B1(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__a21bo_1 _10788_ (.A1(_03355_),
    .A2(_03373_),
    .B1_N(_03372_),
    .X(_03514_));
 sky130_fd_sc_hd__and3_1 _10789_ (.A(_03380_),
    .B(_03412_),
    .C(_03413_),
    .X(_03515_));
 sky130_fd_sc_hd__a21o_1 _10790_ (.A1(_03379_),
    .A2(_03415_),
    .B1(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__or2b_1 _10791_ (.A(_03347_),
    .B_N(_03345_),
    .X(_03517_));
 sky130_fd_sc_hd__nand3_1 _10792_ (.A(_03733_),
    .B(_04251_),
    .C(_03348_),
    .Y(_03519_));
 sky130_fd_sc_hd__a22oi_1 _10793_ (.A1(_06442_),
    .A2(_00093_),
    .B1(_04520_),
    .B2(_06444_),
    .Y(_03520_));
 sky130_fd_sc_hd__and4_1 _10794_ (.A(_00506_),
    .B(_03604_),
    .C(_04445_),
    .D(_00085_),
    .X(_03521_));
 sky130_fd_sc_hd__nor2_1 _10795_ (.A(_03520_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand2_1 _10796_ (.A(_02965_),
    .B(_04380_),
    .Y(_03523_));
 sky130_fd_sc_hd__xnor2_1 _10797_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__buf_2 _10798_ (.A(_06439_),
    .X(_03525_));
 sky130_fd_sc_hd__a31o_1 _10799_ (.A1(_03525_),
    .A2(_04316_),
    .A3(_03343_),
    .B1(_03342_),
    .X(_03526_));
 sky130_fd_sc_hd__xor2_1 _10800_ (.A(_03524_),
    .B(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__and2_1 _10801_ (.A(_03722_),
    .B(_04316_),
    .X(_03528_));
 sky130_fd_sc_hd__xnor2_1 _10802_ (.A(_03527_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__a21oi_1 _10803_ (.A1(_03517_),
    .A2(_03519_),
    .B1(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__and3_1 _10804_ (.A(_03517_),
    .B(_03519_),
    .C(_03529_),
    .X(_03531_));
 sky130_fd_sc_hd__nor2_2 _10805_ (.A(_03530_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2_1 _10806_ (.A(_03798_),
    .B(_04262_),
    .Y(_03533_));
 sky130_fd_sc_hd__xnor2_4 _10807_ (.A(_03532_),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a211oi_1 _10808_ (.A1(_03165_),
    .A2(_03169_),
    .B1(_03368_),
    .C1(_03369_),
    .Y(_03535_));
 sky130_fd_sc_hd__a21o_1 _10809_ (.A1(_03399_),
    .A2(_03408_),
    .B1(_03407_),
    .X(_03536_));
 sky130_fd_sc_hd__o21bai_1 _10810_ (.A1(_03395_),
    .A2(_03398_),
    .B1_N(_03396_),
    .Y(_03537_));
 sky130_fd_sc_hd__a22o_1 _10811_ (.A1(_03443_),
    .A2(_04649_),
    .B1(_00040_),
    .B2(_00281_),
    .X(_03538_));
 sky130_fd_sc_hd__nand4_2 _10812_ (.A(_02983_),
    .B(_02980_),
    .C(_04649_),
    .D(_04714_),
    .Y(_03540_));
 sky130_fd_sc_hd__a22o_1 _10813_ (.A1(_03486_),
    .A2(_04596_),
    .B1(_03538_),
    .B2(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__nand4_2 _10814_ (.A(_02987_),
    .B(_04596_),
    .C(_03538_),
    .D(_03540_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand3_2 _10815_ (.A(_03537_),
    .B(_03541_),
    .C(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__a21o_1 _10816_ (.A1(_03541_),
    .A2(_03542_),
    .B1(_03537_),
    .X(_03544_));
 sky130_fd_sc_hd__nand2_1 _10817_ (.A(_03360_),
    .B(_03362_),
    .Y(_03545_));
 sky130_fd_sc_hd__a21o_1 _10818_ (.A1(_03543_),
    .A2(_03544_),
    .B1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__nand3_1 _10819_ (.A(_03545_),
    .B(_03543_),
    .C(_03544_),
    .Y(_03547_));
 sky130_fd_sc_hd__and3_1 _10820_ (.A(_03536_),
    .B(_03546_),
    .C(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__a21oi_1 _10821_ (.A1(_03546_),
    .A2(_03547_),
    .B1(_03536_),
    .Y(_03549_));
 sky130_fd_sc_hd__a211o_1 _10822_ (.A1(_03363_),
    .A2(_03367_),
    .B1(_03548_),
    .C1(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__o211ai_1 _10823_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03363_),
    .C1(_03367_),
    .Y(_03552_));
 sky130_fd_sc_hd__o211a_1 _10824_ (.A1(_03368_),
    .A2(_03535_),
    .B1(_03551_),
    .C1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a211oi_1 _10825_ (.A1(_03551_),
    .A2(_03552_),
    .B1(_03368_),
    .C1(_03535_),
    .Y(_03554_));
 sky130_fd_sc_hd__nor2_1 _10826_ (.A(_03553_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__xnor2_1 _10827_ (.A(_03534_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__xnor2_1 _10828_ (.A(_03516_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__xor2_2 _10829_ (.A(_03514_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__o21bai_1 _10830_ (.A1(_03419_),
    .A2(_03420_),
    .B1_N(_03421_),
    .Y(_03559_));
 sky130_fd_sc_hd__a22o_1 _10831_ (.A1(_02948_),
    .A2(_06518_),
    .B1(_00412_),
    .B2(_02894_),
    .X(_03560_));
 sky130_fd_sc_hd__nand4_1 _10832_ (.A(_00049_),
    .B(_00046_),
    .C(_05252_),
    .D(_00412_),
    .Y(_03562_));
 sky130_fd_sc_hd__a22o_1 _10833_ (.A1(_03002_),
    .A2(_00002_),
    .B1(_03560_),
    .B2(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__nand4_1 _10834_ (.A(_00058_),
    .B(_00002_),
    .C(_03560_),
    .D(_03562_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand3_1 _10835_ (.A(_03559_),
    .B(_03563_),
    .C(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a21o_1 _10836_ (.A1(_03563_),
    .A2(_03564_),
    .B1(_03559_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_1 _10837_ (.A(_03383_),
    .B(_03385_),
    .Y(_03567_));
 sky130_fd_sc_hd__a21o_1 _10838_ (.A1(_03565_),
    .A2(_03566_),
    .B1(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__nand3_1 _10839_ (.A(_03567_),
    .B(_03565_),
    .C(_03566_),
    .Y(_03569_));
 sky130_fd_sc_hd__a21bo_1 _10840_ (.A1(_03388_),
    .A2(_03387_),
    .B1_N(_03386_),
    .X(_03570_));
 sky130_fd_sc_hd__nand3_4 _10841_ (.A(_03568_),
    .B(_03569_),
    .C(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__a21o_1 _10842_ (.A1(_03568_),
    .A2(_03569_),
    .B1(_03570_),
    .X(_03573_));
 sky130_fd_sc_hd__a22oi_1 _10843_ (.A1(_01146_),
    .A2(_00445_),
    .B1(_00550_),
    .B2(_01147_),
    .Y(_03574_));
 sky130_fd_sc_hd__and4_1 _10844_ (.A(_00124_),
    .B(_00125_),
    .C(_06603_),
    .D(_06605_),
    .X(_03575_));
 sky130_fd_sc_hd__nor2_1 _10845_ (.A(_03574_),
    .B(_03575_),
    .Y(_03576_));
 sky130_fd_sc_hd__nand2_1 _10846_ (.A(_00270_),
    .B(_04789_),
    .Y(_03577_));
 sky130_fd_sc_hd__xnor2_1 _10847_ (.A(_03576_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__a22o_1 _10848_ (.A1(_00096_),
    .A2(_05025_),
    .B1(_06623_),
    .B2(_00095_),
    .X(_03579_));
 sky130_fd_sc_hd__nand4_1 _10849_ (.A(_00086_),
    .B(_00462_),
    .C(_05025_),
    .D(_06623_),
    .Y(_03580_));
 sky130_fd_sc_hd__and2_1 _10850_ (.A(_03152_),
    .B(_06580_),
    .X(_03581_));
 sky130_fd_sc_hd__nand3_1 _10851_ (.A(_03579_),
    .B(_03580_),
    .C(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__a21o_1 _10852_ (.A1(_03579_),
    .A2(_03580_),
    .B1(_03581_),
    .X(_03583_));
 sky130_fd_sc_hd__a21bo_1 _10853_ (.A1(_03403_),
    .A2(_03401_),
    .B1_N(_03402_),
    .X(_03584_));
 sky130_fd_sc_hd__and3_1 _10854_ (.A(_03582_),
    .B(_03583_),
    .C(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _10855_ (.A1(_03582_),
    .A2(_03583_),
    .B1(_03584_),
    .X(_03586_));
 sky130_fd_sc_hd__or2b_1 _10856_ (.A(_03585_),
    .B_N(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__xnor2_1 _10857_ (.A(_03578_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__a21oi_2 _10858_ (.A1(_03571_),
    .A2(_03573_),
    .B1(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__and3_1 _10859_ (.A(_03588_),
    .B(_03571_),
    .C(_03573_),
    .X(_03590_));
 sky130_fd_sc_hd__a211oi_4 _10860_ (.A1(_03437_),
    .A2(_03439_),
    .B1(_03589_),
    .C1(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__o211a_1 _10861_ (.A1(_03589_),
    .A2(_03590_),
    .B1(_03437_),
    .C1(_03439_),
    .X(_03592_));
 sky130_fd_sc_hd__a211oi_4 _10862_ (.A1(_03393_),
    .A2(_03413_),
    .B1(_03591_),
    .C1(_03592_),
    .Y(_03594_));
 sky130_fd_sc_hd__o211a_1 _10863_ (.A1(_03591_),
    .A2(_03592_),
    .B1(_03393_),
    .C1(_03413_),
    .X(_03595_));
 sky130_fd_sc_hd__and3_1 _10864_ (.A(_03460_),
    .B(_03461_),
    .C(_03462_),
    .X(_03596_));
 sky130_fd_sc_hd__and4_1 _10865_ (.A(_03439_),
    .B(_03440_),
    .C(_03463_),
    .D(_03464_),
    .X(_03597_));
 sky130_fd_sc_hd__nand2_1 _10866_ (.A(_03433_),
    .B(_03435_),
    .Y(_03598_));
 sky130_fd_sc_hd__a21bo_1 _10867_ (.A1(_03447_),
    .A2(_03457_),
    .B1_N(_03456_),
    .X(_03599_));
 sky130_fd_sc_hd__a22oi_1 _10868_ (.A1(_06630_),
    .A2(_05445_),
    .B1(_05509_),
    .B2(_06631_),
    .Y(_03600_));
 sky130_fd_sc_hd__and4_1 _10869_ (.A(_06598_),
    .B(_06599_),
    .C(_06489_),
    .D(_05498_),
    .X(_03601_));
 sky130_fd_sc_hd__nor2_1 _10870_ (.A(_03600_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand2_1 _10871_ (.A(net121),
    .B(_06477_),
    .Y(_03603_));
 sky130_fd_sc_hd__xnor2_1 _10872_ (.A(_03602_),
    .B(_03603_),
    .Y(_03605_));
 sky130_fd_sc_hd__a22oi_2 _10873_ (.A1(_02658_),
    .A2(_05638_),
    .B1(_00163_),
    .B2(_02593_),
    .Y(_03606_));
 sky130_fd_sc_hd__and4_1 _10874_ (.A(_06585_),
    .B(_06583_),
    .C(_05638_),
    .D(_06537_),
    .X(_03607_));
 sky130_fd_sc_hd__nand2_1 _10875_ (.A(_02712_),
    .B(_03424_),
    .Y(_03608_));
 sky130_fd_sc_hd__or3_1 _10876_ (.A(_03606_),
    .B(_03607_),
    .C(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__o21ai_1 _10877_ (.A1(_03606_),
    .A2(_03607_),
    .B1(_03608_),
    .Y(_03610_));
 sky130_fd_sc_hd__a21bo_1 _10878_ (.A1(_03428_),
    .A2(_03426_),
    .B1_N(_03427_),
    .X(_03611_));
 sky130_fd_sc_hd__nand3_1 _10879_ (.A(_03609_),
    .B(_03610_),
    .C(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__a21o_1 _10880_ (.A1(_03609_),
    .A2(_03610_),
    .B1(_03611_),
    .X(_03613_));
 sky130_fd_sc_hd__nand3_1 _10881_ (.A(_03605_),
    .B(_03612_),
    .C(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__a21o_1 _10882_ (.A1(_03612_),
    .A2(_03613_),
    .B1(_03605_),
    .X(_03616_));
 sky130_fd_sc_hd__nand3_2 _10883_ (.A(_03599_),
    .B(_03614_),
    .C(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__a21o_1 _10884_ (.A1(_03614_),
    .A2(_03616_),
    .B1(_03599_),
    .X(_03618_));
 sky130_fd_sc_hd__nand3_2 _10885_ (.A(_03598_),
    .B(_03617_),
    .C(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__a21o_1 _10886_ (.A1(_03617_),
    .A2(_03618_),
    .B1(_03598_),
    .X(_03620_));
 sky130_fd_sc_hd__nand2_1 _10887_ (.A(_03451_),
    .B(_03453_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_1 _10888_ (.A(_02528_),
    .B(_03247_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand4_1 _10889_ (.A(_02431_),
    .B(_02229_),
    .C(_00783_),
    .D(_05884_),
    .Y(_03623_));
 sky130_fd_sc_hd__a22o_1 _10890_ (.A1(_02485_),
    .A2(_00785_),
    .B1(_03082_),
    .B2(_06565_),
    .X(_03624_));
 sky130_fd_sc_hd__nand3b_1 _10891_ (.A_N(_03622_),
    .B(_03623_),
    .C(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__a21bo_1 _10892_ (.A1(_03624_),
    .A2(_03623_),
    .B1_N(_03622_),
    .X(_03627_));
 sky130_fd_sc_hd__nand3_1 _10893_ (.A(_03445_),
    .B(_03625_),
    .C(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__a21o_1 _10894_ (.A1(_03625_),
    .A2(_03627_),
    .B1(_03445_),
    .X(_03629_));
 sky130_fd_sc_hd__nand3_1 _10895_ (.A(_03621_),
    .B(_03628_),
    .C(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__a21o_1 _10896_ (.A1(_03628_),
    .A2(_03629_),
    .B1(_03621_),
    .X(_03631_));
 sky130_fd_sc_hd__nand4_2 _10897_ (.A(_02388_),
    .B(_05970_),
    .C(_03630_),
    .D(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__a22o_1 _10898_ (.A1(_02388_),
    .A2(_05970_),
    .B1(_03630_),
    .B2(_03631_),
    .X(_03633_));
 sky130_fd_sc_hd__nand3b_2 _10899_ (.A_N(_03460_),
    .B(_03632_),
    .C(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__a21bo_1 _10900_ (.A1(_03632_),
    .A2(_03633_),
    .B1_N(_03460_),
    .X(_03635_));
 sky130_fd_sc_hd__a22o_1 _10901_ (.A1(_03619_),
    .A2(_03620_),
    .B1(_03634_),
    .B2(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__nand4_2 _10902_ (.A(_03619_),
    .B(_03620_),
    .C(_03634_),
    .D(_03635_),
    .Y(_03638_));
 sky130_fd_sc_hd__o211a_1 _10903_ (.A1(_03596_),
    .A2(_03597_),
    .B1(_03636_),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a211oi_1 _10904_ (.A1(_03636_),
    .A2(_03638_),
    .B1(_03596_),
    .C1(_03597_),
    .Y(_03640_));
 sky130_fd_sc_hd__nor4_1 _10905_ (.A(_03594_),
    .B(_03595_),
    .C(_03639_),
    .D(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__o22a_1 _10906_ (.A1(_03594_),
    .A2(_03595_),
    .B1(_03639_),
    .B2(_03640_),
    .X(_03642_));
 sky130_fd_sc_hd__nor2_1 _10907_ (.A(_03641_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__and2b_1 _10908_ (.A_N(_03469_),
    .B(_03467_),
    .X(_03644_));
 sky130_fd_sc_hd__a21oi_1 _10909_ (.A1(_03416_),
    .A2(_03470_),
    .B1(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__xnor2_2 _10910_ (.A(_03643_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__xnor2_2 _10911_ (.A(_03558_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__and2b_1 _10912_ (.A_N(_03473_),
    .B(_03471_),
    .X(_03648_));
 sky130_fd_sc_hd__a21oi_2 _10913_ (.A1(_03377_),
    .A2(_03474_),
    .B1(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__xnor2_2 _10914_ (.A(_03647_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__xnor2_4 _10915_ (.A(_03513_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__inv_2 _10916_ (.A(_03334_),
    .Y(_03652_));
 sky130_fd_sc_hd__or2_1 _10917_ (.A(_03475_),
    .B(_03477_),
    .X(_03653_));
 sky130_fd_sc_hd__o21ai_4 _10918_ (.A1(_03652_),
    .A2(_03478_),
    .B1(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__xor2_4 _10919_ (.A(_03651_),
    .B(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__xnor2_1 _10920_ (.A(_03511_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__a21o_1 _10921_ (.A1(_03509_),
    .A2(_03510_),
    .B1(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__nand3_1 _10922_ (.A(_03509_),
    .B(_03510_),
    .C(_03656_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(_03657_),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__nor2_1 _10924_ (.A(_03294_),
    .B(_03485_),
    .Y(_03661_));
 sky130_fd_sc_hd__nand2_1 _10925_ (.A(_03331_),
    .B(_03484_),
    .Y(_03662_));
 sky130_fd_sc_hd__nor2_1 _10926_ (.A(_03331_),
    .B(_03484_),
    .Y(_03663_));
 sky130_fd_sc_hd__a221o_1 _10927_ (.A1(_03328_),
    .A2(_03662_),
    .B1(_03661_),
    .B2(_03296_),
    .C1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__a31oi_1 _10928_ (.A1(_02703_),
    .A2(_03295_),
    .A3(_03661_),
    .B1(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _10929_ (.A(_03660_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(_03660_),
    .B(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__o21ai_1 _10931_ (.A1(_02544_),
    .A2(_02554_),
    .B1(_02563_),
    .Y(_03668_));
 sky130_fd_sc_hd__and3b_1 _10932_ (.A_N(_02564_),
    .B(_03314_),
    .C(_03668_),
    .X(_03670_));
 sky130_fd_sc_hd__a21o_1 _10933_ (.A1(_03318_),
    .A2(_03490_),
    .B1(_02351_),
    .X(_03671_));
 sky130_fd_sc_hd__or2_1 _10934_ (.A(_02764_),
    .B(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__nand2_1 _10935_ (.A(_02764_),
    .B(_03671_),
    .Y(_03673_));
 sky130_fd_sc_hd__a2bb2o_1 _10936_ (.A1_N(_04197_),
    .A2_N(_02941_),
    .B1(_02731_),
    .B2(\AuI.result[4] ),
    .X(_03674_));
 sky130_fd_sc_hd__clkbuf_4 _10937_ (.A(_02718_),
    .X(_03675_));
 sky130_fd_sc_hd__a22o_1 _10938_ (.A1(_02350_),
    .A2(_02742_),
    .B1(_02943_),
    .B2(_04133_),
    .X(_03676_));
 sky130_fd_sc_hd__a221o_1 _10939_ (.A1(\MuI.result[4] ),
    .A2(_02736_),
    .B1(_02707_),
    .B2(_02764_),
    .C1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__a221o_1 _10940_ (.A1(_04262_),
    .A2(_03675_),
    .B1(_02721_),
    .B2(_02345_),
    .C1(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__a211o_1 _10941_ (.A1(\FuI.Integer[4] ),
    .A2(_06056_),
    .B1(_03674_),
    .C1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__a31o_1 _10942_ (.A1(_03489_),
    .A2(_03672_),
    .A3(_03673_),
    .B1(_03679_),
    .X(_03681_));
 sky130_fd_sc_hd__a311o_1 _10943_ (.A1(_03134_),
    .A2(_03666_),
    .A3(_03667_),
    .B1(_03670_),
    .C1(_03681_),
    .X(_03682_));
 sky130_fd_sc_hd__a31o_2 _10944_ (.A1(_02752_),
    .A2(_03506_),
    .A3(_03508_),
    .B1(_03682_),
    .X(net95));
 sky130_fd_sc_hd__or2b_1 _10945_ (.A(_02345_),
    .B_N(_04197_),
    .X(_03683_));
 sky130_fd_sc_hd__and2b_1 _10946_ (.A_N(_02883_),
    .B(_03322_),
    .X(_03684_));
 sky130_fd_sc_hd__a2111o_1 _10947_ (.A1(_02769_),
    .A2(_03321_),
    .B1(_03684_),
    .C1(_03317_),
    .D1(_02762_),
    .X(_03685_));
 sky130_fd_sc_hd__nand2_1 _10948_ (.A(_03683_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__o21a_1 _10949_ (.A1(_02764_),
    .A2(_03503_),
    .B1(_03683_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(_03686_),
    .A1(_03687_),
    .S(_02928_),
    .X(_03688_));
 sky130_fd_sc_hd__xnor2_1 _10951_ (.A(_02760_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _10952_ (.A(_03657_),
    .B(_03667_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand2_2 _10953_ (.A(_03651_),
    .B(_03654_),
    .Y(_03692_));
 sky130_fd_sc_hd__nand2_1 _10954_ (.A(_03511_),
    .B(_03655_),
    .Y(_03693_));
 sky130_fd_sc_hd__a31o_1 _10955_ (.A1(_03820_),
    .A2(_04262_),
    .A3(_03532_),
    .B1(_03530_),
    .X(_03694_));
 sky130_fd_sc_hd__and2b_1 _10956_ (.A_N(_03556_),
    .B(_03516_),
    .X(_03695_));
 sky130_fd_sc_hd__a21o_2 _10957_ (.A1(_03514_),
    .A2(_03557_),
    .B1(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__and2_1 _10958_ (.A(_03534_),
    .B(_03555_),
    .X(_03697_));
 sky130_fd_sc_hd__and3_1 _10959_ (.A(_03539_),
    .B(_00678_),
    .C(_00085_),
    .X(_03698_));
 sky130_fd_sc_hd__a22o_1 _10960_ (.A1(_00678_),
    .A2(_00085_),
    .B1(_00047_),
    .B2(_03539_),
    .X(_03699_));
 sky130_fd_sc_hd__a21bo_1 _10961_ (.A1(_04596_),
    .A2(_03698_),
    .B1_N(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(_03658_),
    .B(_04456_),
    .Y(_03702_));
 sky130_fd_sc_hd__xor2_4 _10963_ (.A(_03700_),
    .B(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__a31o_2 _10964_ (.A1(_03525_),
    .A2(_04380_),
    .A3(_03522_),
    .B1(_03521_),
    .X(_03704_));
 sky130_fd_sc_hd__xor2_4 _10965_ (.A(_03703_),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__nand2_1 _10966_ (.A(net60),
    .B(_04380_),
    .Y(_03706_));
 sky130_fd_sc_hd__clkinv_2 _10967_ (.A(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__xnor2_4 _10968_ (.A(_03705_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__and2_1 _10969_ (.A(_03524_),
    .B(_03526_),
    .X(_03709_));
 sky130_fd_sc_hd__a21o_1 _10970_ (.A1(_03527_),
    .A2(_03528_),
    .B1(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_4 _10971_ (.A(_03708_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__nand2_1 _10972_ (.A(_00502_),
    .B(_04316_),
    .Y(_03712_));
 sky130_fd_sc_hd__xnor2_4 _10973_ (.A(_03711_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__a211oi_1 _10974_ (.A1(_03363_),
    .A2(_03367_),
    .B1(_03548_),
    .C1(_03549_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21o_1 _10975_ (.A1(_03578_),
    .A2(_03586_),
    .B1(_03585_),
    .X(_03715_));
 sky130_fd_sc_hd__o21bai_1 _10976_ (.A1(_03574_),
    .A2(_03577_),
    .B1_N(_03575_),
    .Y(_03716_));
 sky130_fd_sc_hd__a22o_1 _10977_ (.A1(_00289_),
    .A2(_00033_),
    .B1(_06612_),
    .B2(_00290_),
    .X(_03717_));
 sky130_fd_sc_hd__nand4_1 _10978_ (.A(_00281_),
    .B(_03443_),
    .C(_00040_),
    .D(_04789_),
    .Y(_03718_));
 sky130_fd_sc_hd__a22o_1 _10979_ (.A1(_03486_),
    .A2(_00059_),
    .B1(_03717_),
    .B2(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__nand4_1 _10980_ (.A(_00345_),
    .B(_00059_),
    .C(_03717_),
    .D(_03718_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand3_2 _10981_ (.A(_03716_),
    .B(_03719_),
    .C(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__a21o_1 _10982_ (.A1(_03719_),
    .A2(_03720_),
    .B1(_03716_),
    .X(_03723_));
 sky130_fd_sc_hd__nand2_1 _10983_ (.A(_03540_),
    .B(_03542_),
    .Y(_03724_));
 sky130_fd_sc_hd__a21o_1 _10984_ (.A1(_03721_),
    .A2(_03723_),
    .B1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__nand3_2 _10985_ (.A(_03724_),
    .B(_03721_),
    .C(_03723_),
    .Y(_03726_));
 sky130_fd_sc_hd__and3_1 _10986_ (.A(_03715_),
    .B(_03725_),
    .C(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__a21oi_1 _10987_ (.A1(_03725_),
    .A2(_03726_),
    .B1(_03715_),
    .Y(_03728_));
 sky130_fd_sc_hd__a211o_1 _10988_ (.A1(_03543_),
    .A2(_03547_),
    .B1(_03727_),
    .C1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__o211ai_1 _10989_ (.A1(_03727_),
    .A2(_03728_),
    .B1(_03543_),
    .C1(_03547_),
    .Y(_03730_));
 sky130_fd_sc_hd__o211ai_2 _10990_ (.A1(_03548_),
    .A2(_03714_),
    .B1(_03729_),
    .C1(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__a211o_1 _10991_ (.A1(_03729_),
    .A2(_03730_),
    .B1(_03548_),
    .C1(_03714_),
    .X(_03732_));
 sky130_fd_sc_hd__nand3_1 _10992_ (.A(_03713_),
    .B(_03731_),
    .C(_03732_),
    .Y(_03734_));
 sky130_fd_sc_hd__a21o_1 _10993_ (.A1(_03731_),
    .A2(_03732_),
    .B1(_03713_),
    .X(_03735_));
 sky130_fd_sc_hd__o211ai_1 _10994_ (.A1(_03591_),
    .A2(_03594_),
    .B1(_03734_),
    .C1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__a211o_1 _10995_ (.A1(_03734_),
    .A2(_03735_),
    .B1(_03591_),
    .C1(_03594_),
    .X(_03737_));
 sky130_fd_sc_hd__o211a_1 _10996_ (.A1(_03553_),
    .A2(_03697_),
    .B1(_03736_),
    .C1(_03737_),
    .X(_03738_));
 sky130_fd_sc_hd__a211oi_1 _10997_ (.A1(_03736_),
    .A2(_03737_),
    .B1(_03553_),
    .C1(_03697_),
    .Y(_03739_));
 sky130_fd_sc_hd__or2_1 _10998_ (.A(_03738_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__nand3_2 _10999_ (.A(_03588_),
    .B(_03571_),
    .C(_03573_),
    .Y(_03741_));
 sky130_fd_sc_hd__o21bai_1 _11000_ (.A1(_03600_),
    .A2(_03603_),
    .B1_N(_03601_),
    .Y(_03742_));
 sky130_fd_sc_hd__a22o_1 _11001_ (.A1(_02948_),
    .A2(_06562_),
    .B1(_06476_),
    .B2(_00028_),
    .X(_03743_));
 sky130_fd_sc_hd__nand4_1 _11002_ (.A(_02894_),
    .B(_00046_),
    .C(_00412_),
    .D(_00530_),
    .Y(_03745_));
 sky130_fd_sc_hd__a22o_1 _11003_ (.A1(_03002_),
    .A2(_06561_),
    .B1(_03743_),
    .B2(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__nand4_1 _11004_ (.A(_00058_),
    .B(_06561_),
    .C(_03743_),
    .D(_03745_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand3_1 _11005_ (.A(_03742_),
    .B(_03746_),
    .C(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__a21o_1 _11006_ (.A1(_03746_),
    .A2(_03747_),
    .B1(_03742_),
    .X(_03749_));
 sky130_fd_sc_hd__nand2_1 _11007_ (.A(_03562_),
    .B(_03564_),
    .Y(_03750_));
 sky130_fd_sc_hd__a21o_1 _11008_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_03750_),
    .X(_03751_));
 sky130_fd_sc_hd__nand3_2 _11009_ (.A(_03750_),
    .B(_03748_),
    .C(_03749_),
    .Y(_03752_));
 sky130_fd_sc_hd__a21bo_1 _11010_ (.A1(_03567_),
    .A2(_03566_),
    .B1_N(_03565_),
    .X(_03753_));
 sky130_fd_sc_hd__nand3_4 _11011_ (.A(_03751_),
    .B(_03752_),
    .C(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__a21o_1 _11012_ (.A1(_03751_),
    .A2(_03752_),
    .B1(_03753_),
    .X(_03756_));
 sky130_fd_sc_hd__a22oi_1 _11013_ (.A1(_01146_),
    .A2(_00550_),
    .B1(_00197_),
    .B2(_01147_),
    .Y(_03757_));
 sky130_fd_sc_hd__and4_1 _11014_ (.A(_00124_),
    .B(_00125_),
    .C(_06605_),
    .D(_06591_),
    .X(_03758_));
 sky130_fd_sc_hd__nor2_1 _11015_ (.A(_03757_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand2_1 _11016_ (.A(_03324_),
    .B(_00445_),
    .Y(_03760_));
 sky130_fd_sc_hd__xnor2_2 _11017_ (.A(_03759_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__a22o_1 _11018_ (.A1(_00096_),
    .A2(_05101_),
    .B1(_06517_),
    .B2(_00095_),
    .X(_03762_));
 sky130_fd_sc_hd__nand4_1 _11019_ (.A(_00086_),
    .B(_00081_),
    .C(_06623_),
    .D(_06517_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand4_1 _11020_ (.A(_00262_),
    .B(_00421_),
    .C(_03762_),
    .D(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__a22o_1 _11021_ (.A1(_00088_),
    .A2(_05036_),
    .B1(_03762_),
    .B2(_03763_),
    .X(_03765_));
 sky130_fd_sc_hd__a21bo_1 _11022_ (.A1(_03579_),
    .A2(_03581_),
    .B1_N(_03580_),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _11023_ (.A(_03764_),
    .B(_03765_),
    .C(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__a21o_1 _11024_ (.A1(_03764_),
    .A2(_03765_),
    .B1(_03767_),
    .X(_03769_));
 sky130_fd_sc_hd__and2b_1 _11025_ (.A_N(_03768_),
    .B(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__xor2_2 _11026_ (.A(_03761_),
    .B(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__a21oi_2 _11027_ (.A1(_03754_),
    .A2(_03756_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__and3_1 _11028_ (.A(_03771_),
    .B(_03754_),
    .C(_03756_),
    .X(_03773_));
 sky130_fd_sc_hd__a211oi_4 _11029_ (.A1(_03617_),
    .A2(_03619_),
    .B1(_03772_),
    .C1(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__o211a_1 _11030_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03617_),
    .C1(_03619_),
    .X(_03775_));
 sky130_fd_sc_hd__a211oi_4 _11031_ (.A1(_03571_),
    .A2(_03741_),
    .B1(_03774_),
    .C1(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__o211a_1 _11032_ (.A1(_03774_),
    .A2(_03775_),
    .B1(_03571_),
    .C1(_03741_),
    .X(_03778_));
 sky130_fd_sc_hd__nand2_1 _11033_ (.A(_03612_),
    .B(_03614_),
    .Y(_03779_));
 sky130_fd_sc_hd__a21bo_1 _11034_ (.A1(_03621_),
    .A2(_03629_),
    .B1_N(_03628_),
    .X(_03780_));
 sky130_fd_sc_hd__a22oi_1 _11035_ (.A1(_00011_),
    .A2(_05509_),
    .B1(_05574_),
    .B2(_00012_),
    .Y(_03781_));
 sky130_fd_sc_hd__and4_1 _11036_ (.A(_02754_),
    .B(_02797_),
    .C(_00398_),
    .D(_03424_),
    .X(_03782_));
 sky130_fd_sc_hd__nor2_1 _11037_ (.A(_03781_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(_06608_),
    .B(_06546_),
    .Y(_03784_));
 sky130_fd_sc_hd__xnor2_1 _11039_ (.A(_03783_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__a22oi_2 _11040_ (.A1(_06583_),
    .A2(_06537_),
    .B1(_05756_),
    .B2(_06585_),
    .Y(_03786_));
 sky130_fd_sc_hd__and4_1 _11041_ (.A(_00414_),
    .B(_06622_),
    .C(net130),
    .D(net129),
    .X(_03787_));
 sky130_fd_sc_hd__nand2_1 _11042_ (.A(_06680_),
    .B(_00382_),
    .Y(_03788_));
 sky130_fd_sc_hd__or3_1 _11043_ (.A(_03786_),
    .B(_03787_),
    .C(_03788_),
    .X(_03789_));
 sky130_fd_sc_hd__o21ai_1 _11044_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_03788_),
    .Y(_03790_));
 sky130_fd_sc_hd__o21bai_1 _11045_ (.A1(_03606_),
    .A2(_03608_),
    .B1_N(_03607_),
    .Y(_03791_));
 sky130_fd_sc_hd__nand3_1 _11046_ (.A(_03789_),
    .B(_03790_),
    .C(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__a21o_1 _11047_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03791_),
    .X(_03793_));
 sky130_fd_sc_hd__nand3_1 _11048_ (.A(_03785_),
    .B(_03792_),
    .C(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__a21o_1 _11049_ (.A1(_03792_),
    .A2(_03793_),
    .B1(_03785_),
    .X(_03795_));
 sky130_fd_sc_hd__nand3_2 _11050_ (.A(_03780_),
    .B(_03794_),
    .C(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__a21o_1 _11051_ (.A1(_03794_),
    .A2(_03795_),
    .B1(_03780_),
    .X(_03797_));
 sky130_fd_sc_hd__nand3_2 _11052_ (.A(_03779_),
    .B(_03796_),
    .C(_03797_),
    .Y(_03799_));
 sky130_fd_sc_hd__a21o_1 _11053_ (.A1(_03796_),
    .A2(_03797_),
    .B1(_03779_),
    .X(_03800_));
 sky130_fd_sc_hd__and3_1 _11054_ (.A(_06565_),
    .B(_03082_),
    .C(_00789_),
    .X(_03801_));
 sky130_fd_sc_hd__a22o_1 _11055_ (.A1(_02485_),
    .A2(_03082_),
    .B1(_00789_),
    .B2(_06565_),
    .X(_03802_));
 sky130_fd_sc_hd__a21bo_1 _11056_ (.A1(_02496_),
    .A2(_03801_),
    .B1_N(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__nand2_1 _11057_ (.A(_02539_),
    .B(_03257_),
    .Y(_03804_));
 sky130_fd_sc_hd__xor2_2 _11058_ (.A(_03803_),
    .B(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_03623_),
    .B(_03625_),
    .Y(_03806_));
 sky130_fd_sc_hd__xnor2_1 _11060_ (.A(_03805_),
    .B(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__xor2_1 _11061_ (.A(_03632_),
    .B(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__a21oi_1 _11062_ (.A1(_03799_),
    .A2(_03800_),
    .B1(_03808_),
    .Y(_03810_));
 sky130_fd_sc_hd__and3_1 _11063_ (.A(_03808_),
    .B(_03799_),
    .C(_03800_),
    .X(_03811_));
 sky130_fd_sc_hd__a211o_1 _11064_ (.A1(_03634_),
    .A2(_03638_),
    .B1(_03810_),
    .C1(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__o211ai_1 _11065_ (.A1(_03810_),
    .A2(_03811_),
    .B1(_03634_),
    .C1(_03638_),
    .Y(_03813_));
 sky130_fd_sc_hd__a2bb2o_1 _11066_ (.A1_N(_03776_),
    .A2_N(_03778_),
    .B1(_03812_),
    .B2(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__or4bb_2 _11067_ (.A(_03776_),
    .B(_03778_),
    .C_N(_03812_),
    .D_N(_03813_),
    .X(_03815_));
 sky130_fd_sc_hd__o211a_1 _11068_ (.A1(_03639_),
    .A2(_03641_),
    .B1(_03814_),
    .C1(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__a211o_1 _11069_ (.A1(_03814_),
    .A2(_03815_),
    .B1(_03639_),
    .C1(_03641_),
    .X(_03817_));
 sky130_fd_sc_hd__and2b_1 _11070_ (.A_N(_03816_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__xnor2_2 _11071_ (.A(_03740_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__and2b_1 _11072_ (.A_N(_03645_),
    .B(_03643_),
    .X(_03821_));
 sky130_fd_sc_hd__a21oi_2 _11073_ (.A1(_03558_),
    .A2(_03646_),
    .B1(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__xnor2_4 _11074_ (.A(_03819_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__xor2_4 _11075_ (.A(_03696_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_1 _11076_ (.A(_03647_),
    .B(_03649_),
    .Y(_03825_));
 sky130_fd_sc_hd__nor2_1 _11077_ (.A(_03647_),
    .B(_03649_),
    .Y(_03826_));
 sky130_fd_sc_hd__a21oi_2 _11078_ (.A1(_03513_),
    .A2(_03825_),
    .B1(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__xnor2_4 _11079_ (.A(_03824_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _11080_ (.A(_03694_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__a21oi_1 _11081_ (.A1(_03692_),
    .A2(_03693_),
    .B1(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__and3_1 _11082_ (.A(_03692_),
    .B(_03693_),
    .C(_03829_),
    .X(_03832_));
 sky130_fd_sc_hd__nor2_1 _11083_ (.A(_03830_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__a21oi_1 _11084_ (.A1(_03691_),
    .A2(_03833_),
    .B1(_06428_),
    .Y(_03834_));
 sky130_fd_sc_hd__o21a_1 _11085_ (.A1(_03691_),
    .A2(_03833_),
    .B1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__nor3_1 _11086_ (.A(_02530_),
    .B(_02544_),
    .C(_02564_),
    .Y(_03836_));
 sky130_fd_sc_hd__nor2_1 _11087_ (.A(_02565_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__a21oi_1 _11088_ (.A1(_02764_),
    .A2(_03671_),
    .B1(_02350_),
    .Y(_03838_));
 sky130_fd_sc_hd__a21oi_1 _11089_ (.A1(_02760_),
    .A2(_03838_),
    .B1(_02711_),
    .Y(_03839_));
 sky130_fd_sc_hd__o21a_1 _11090_ (.A1(_02760_),
    .A2(_03838_),
    .B1(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a2bb2o_1 _11091_ (.A1_N(_03306_),
    .A2_N(_02760_),
    .B1(_02722_),
    .B2(_02388_),
    .X(_03841_));
 sky130_fd_sc_hd__a2bb2o_1 _11092_ (.A1_N(_04262_),
    .A2_N(_02728_),
    .B1(_03675_),
    .B2(_04327_),
    .X(_03843_));
 sky130_fd_sc_hd__and3_1 _11093_ (.A(_02388_),
    .B(_04262_),
    .C(_02743_),
    .X(_03844_));
 sky130_fd_sc_hd__a221o_1 _11094_ (.A1(\MuI.result[5] ),
    .A2(_02737_),
    .B1(_02945_),
    .B2(_04197_),
    .C1(_03844_),
    .X(_03845_));
 sky130_fd_sc_hd__a221o_1 _11095_ (.A1(\FuI.Integer[5] ),
    .A2(_02931_),
    .B1(_02938_),
    .B2(\AuI.result[5] ),
    .C1(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__or4_1 _11096_ (.A(_03840_),
    .B(_03841_),
    .C(_03843_),
    .D(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__a31o_1 _11097_ (.A1(_02552_),
    .A2(_03315_),
    .A3(_03837_),
    .B1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__a211o_2 _11098_ (.A1(_02751_),
    .A2(_03689_),
    .B1(_03835_),
    .C1(_03848_),
    .X(net96));
 sky130_fd_sc_hd__a21o_1 _11099_ (.A1(_02545_),
    .A2(_02553_),
    .B1(_02565_),
    .X(_03849_));
 sky130_fd_sc_hd__a21oi_1 _11100_ (.A1(_03683_),
    .A2(_03685_),
    .B1(_02758_),
    .Y(_03850_));
 sky130_fd_sc_hd__nor2_1 _11101_ (.A(_02759_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__and2_1 _11102_ (.A(_02879_),
    .B(_02886_),
    .X(_03853_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(_03851_),
    .A1(_03853_),
    .S(_02925_),
    .X(_03854_));
 sky130_fd_sc_hd__nand2_1 _11104_ (.A(_02757_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__or2_1 _11105_ (.A(_02757_),
    .B(_03854_),
    .X(_03856_));
 sky130_fd_sc_hd__and2b_1 _11106_ (.A_N(_03708_),
    .B(_03710_),
    .X(_03857_));
 sky130_fd_sc_hd__a31o_1 _11107_ (.A1(_03809_),
    .A2(_04327_),
    .A3(_03711_),
    .B1(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__inv_2 _11108_ (.A(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__o211a_1 _11109_ (.A1(_03591_),
    .A2(_03594_),
    .B1(_03734_),
    .C1(_03735_),
    .X(_03860_));
 sky130_fd_sc_hd__or2_2 _11110_ (.A(_03860_),
    .B(_03738_),
    .X(_03861_));
 sky130_fd_sc_hd__nor4b_1 _11111_ (.A(_03738_),
    .B(_03739_),
    .C(_03816_),
    .D_N(_03817_),
    .Y(_03862_));
 sky130_fd_sc_hd__inv_2 _11112_ (.A(_03731_),
    .Y(_03863_));
 sky130_fd_sc_hd__and3_1 _11113_ (.A(_03713_),
    .B(_03731_),
    .C(_03732_),
    .X(_03864_));
 sky130_fd_sc_hd__and3_1 _11114_ (.A(_03539_),
    .B(_00678_),
    .C(_00047_),
    .X(_03865_));
 sky130_fd_sc_hd__a22o_1 _11115_ (.A1(_00678_),
    .A2(_00047_),
    .B1(_00048_),
    .B2(_06434_),
    .X(_03866_));
 sky130_fd_sc_hd__a21bo_1 _11116_ (.A1(_00059_),
    .A2(_03865_),
    .B1_N(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__nand2_1 _11117_ (.A(_03658_),
    .B(_04531_),
    .Y(_03868_));
 sky130_fd_sc_hd__xor2_4 _11118_ (.A(_03867_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__a32o_2 _11119_ (.A1(_03525_),
    .A2(_04456_),
    .A3(_03699_),
    .B1(_03698_),
    .B2(_04596_),
    .X(_03870_));
 sky130_fd_sc_hd__xor2_4 _11120_ (.A(_03869_),
    .B(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__and2_2 _11121_ (.A(_03722_),
    .B(_04456_),
    .X(_03872_));
 sky130_fd_sc_hd__xnor2_4 _11122_ (.A(_03871_),
    .B(_03872_),
    .Y(_03874_));
 sky130_fd_sc_hd__and2_1 _11123_ (.A(_03703_),
    .B(_03704_),
    .X(_03875_));
 sky130_fd_sc_hd__a21oi_4 _11124_ (.A1(_03705_),
    .A2(_03707_),
    .B1(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__xor2_4 _11125_ (.A(_03874_),
    .B(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(_00502_),
    .B(_04380_),
    .Y(_03878_));
 sky130_fd_sc_hd__xnor2_4 _11127_ (.A(_03877_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__a211oi_1 _11128_ (.A1(_03543_),
    .A2(_03547_),
    .B1(_03727_),
    .C1(_03728_),
    .Y(_03880_));
 sky130_fd_sc_hd__a21o_1 _11129_ (.A1(_03761_),
    .A2(_03769_),
    .B1(_03768_),
    .X(_03881_));
 sky130_fd_sc_hd__o21bai_1 _11130_ (.A1(_03757_),
    .A2(_03760_),
    .B1_N(_03758_),
    .Y(_03882_));
 sky130_fd_sc_hd__a22o_1 _11131_ (.A1(_03443_),
    .A2(_06612_),
    .B1(_04843_),
    .B2(_00290_),
    .X(_03883_));
 sky130_fd_sc_hd__nand4_2 _11132_ (.A(_02983_),
    .B(_02980_),
    .C(_04789_),
    .D(_00445_),
    .Y(_03885_));
 sky130_fd_sc_hd__a22o_1 _11133_ (.A1(_03486_),
    .A2(_04725_),
    .B1(_03883_),
    .B2(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__nand4_2 _11134_ (.A(_00345_),
    .B(_04725_),
    .C(_03883_),
    .D(_03885_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand3_2 _11135_ (.A(_03882_),
    .B(_03886_),
    .C(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__a21o_1 _11136_ (.A1(_03886_),
    .A2(_03887_),
    .B1(_03882_),
    .X(_03889_));
 sky130_fd_sc_hd__nand2_1 _11137_ (.A(_03718_),
    .B(_03720_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _11138_ (.A1(_03888_),
    .A2(_03889_),
    .B1(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__nand3_2 _11139_ (.A(_03890_),
    .B(_03888_),
    .C(_03889_),
    .Y(_03892_));
 sky130_fd_sc_hd__and3_2 _11140_ (.A(_03881_),
    .B(_03891_),
    .C(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__a21oi_1 _11141_ (.A1(_03891_),
    .A2(_03892_),
    .B1(_03881_),
    .Y(_03894_));
 sky130_fd_sc_hd__a211o_1 _11142_ (.A1(_03721_),
    .A2(_03726_),
    .B1(_03893_),
    .C1(_03894_),
    .X(_03896_));
 sky130_fd_sc_hd__o211ai_1 _11143_ (.A1(_03893_),
    .A2(_03894_),
    .B1(_03721_),
    .C1(_03726_),
    .Y(_03897_));
 sky130_fd_sc_hd__o211ai_2 _11144_ (.A1(_03727_),
    .A2(_03880_),
    .B1(_03896_),
    .C1(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__a211o_1 _11145_ (.A1(_03896_),
    .A2(_03897_),
    .B1(_03727_),
    .C1(_03880_),
    .X(_03899_));
 sky130_fd_sc_hd__nand3_1 _11146_ (.A(_03879_),
    .B(_03898_),
    .C(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__a21o_1 _11147_ (.A1(_03898_),
    .A2(_03899_),
    .B1(_03879_),
    .X(_03901_));
 sky130_fd_sc_hd__o211ai_4 _11148_ (.A1(_03774_),
    .A2(_03776_),
    .B1(_03900_),
    .C1(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__a211o_1 _11149_ (.A1(_03900_),
    .A2(_03901_),
    .B1(_03774_),
    .C1(_03776_),
    .X(_03903_));
 sky130_fd_sc_hd__o211ai_4 _11150_ (.A1(_03863_),
    .A2(_03864_),
    .B1(_03902_),
    .C1(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__a211o_1 _11151_ (.A1(_03902_),
    .A2(_03903_),
    .B1(_03863_),
    .C1(_03864_),
    .X(_03905_));
 sky130_fd_sc_hd__or2_1 _11152_ (.A(_03632_),
    .B(_03807_),
    .X(_03907_));
 sky130_fd_sc_hd__nand3_1 _11153_ (.A(_03808_),
    .B(_03799_),
    .C(_03800_),
    .Y(_03908_));
 sky130_fd_sc_hd__nand2_1 _11154_ (.A(_02496_),
    .B(_05895_),
    .Y(_03909_));
 sky130_fd_sc_hd__nand2_1 _11155_ (.A(_02539_),
    .B(_05959_),
    .Y(_03910_));
 sky130_fd_sc_hd__a22o_1 _11156_ (.A1(_02539_),
    .A2(_05895_),
    .B1(_05959_),
    .B2(_02496_),
    .X(_03911_));
 sky130_fd_sc_hd__o21a_1 _11157_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__and2_1 _11158_ (.A(_02229_),
    .B(_05884_),
    .X(_03913_));
 sky130_fd_sc_hd__and3_1 _11159_ (.A(_02442_),
    .B(_05948_),
    .C(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__a31o_1 _11160_ (.A1(_02550_),
    .A2(_05831_),
    .A3(_03802_),
    .B1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__and2_1 _11161_ (.A(_03912_),
    .B(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__nor2_1 _11162_ (.A(_03912_),
    .B(_03915_),
    .Y(_03918_));
 sky130_fd_sc_hd__nor2_1 _11163_ (.A(_03916_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _11164_ (.A(_03792_),
    .B(_03794_),
    .Y(_03920_));
 sky130_fd_sc_hd__and2_1 _11165_ (.A(_03805_),
    .B(_03806_),
    .X(_03921_));
 sky130_fd_sc_hd__a22oi_1 _11166_ (.A1(_00878_),
    .A2(_05574_),
    .B1(_05649_),
    .B2(_00877_),
    .Y(_03922_));
 sky130_fd_sc_hd__and4_1 _11167_ (.A(_02754_),
    .B(_02797_),
    .C(_03424_),
    .D(_00382_),
    .X(_03923_));
 sky130_fd_sc_hd__nor2_1 _11168_ (.A(_03922_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _11169_ (.A(_06608_),
    .B(_03051_),
    .Y(_03925_));
 sky130_fd_sc_hd__xnor2_1 _11170_ (.A(_03924_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__a22oi_2 _11171_ (.A1(_02658_),
    .A2(_00385_),
    .B1(_00783_),
    .B2(_02593_),
    .Y(_03927_));
 sky130_fd_sc_hd__and4_1 _11172_ (.A(_00414_),
    .B(_06622_),
    .C(_05756_),
    .D(_00785_),
    .X(_03929_));
 sky130_fd_sc_hd__nand2_1 _11173_ (.A(_06680_),
    .B(_00163_),
    .Y(_03930_));
 sky130_fd_sc_hd__or3_1 _11174_ (.A(_03927_),
    .B(_03929_),
    .C(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__o21ai_1 _11175_ (.A1(_03927_),
    .A2(_03929_),
    .B1(_03930_),
    .Y(_03932_));
 sky130_fd_sc_hd__o21bai_1 _11176_ (.A1(_03786_),
    .A2(_03788_),
    .B1_N(_03787_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand3_1 _11177_ (.A(_03931_),
    .B(_03932_),
    .C(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__a21o_1 _11178_ (.A1(_03931_),
    .A2(_03932_),
    .B1(_03933_),
    .X(_03935_));
 sky130_fd_sc_hd__nand3_1 _11179_ (.A(_03926_),
    .B(_03934_),
    .C(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__a21o_1 _11180_ (.A1(_03934_),
    .A2(_03935_),
    .B1(_03926_),
    .X(_03937_));
 sky130_fd_sc_hd__nand3_2 _11181_ (.A(_03921_),
    .B(_03936_),
    .C(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hd__a21o_1 _11182_ (.A1(_03936_),
    .A2(_03937_),
    .B1(_03921_),
    .X(_03940_));
 sky130_fd_sc_hd__nand3_2 _11183_ (.A(_03920_),
    .B(_03938_),
    .C(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21o_1 _11184_ (.A1(_03938_),
    .A2(_03940_),
    .B1(_03920_),
    .X(_03942_));
 sky130_fd_sc_hd__and3_1 _11185_ (.A(_03919_),
    .B(_03941_),
    .C(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__a21oi_1 _11186_ (.A1(_03941_),
    .A2(_03942_),
    .B1(_03919_),
    .Y(_03944_));
 sky130_fd_sc_hd__a211oi_2 _11187_ (.A1(_03907_),
    .A2(_03908_),
    .B1(_03943_),
    .C1(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__o211a_1 _11188_ (.A1(_03943_),
    .A2(_03944_),
    .B1(_03907_),
    .C1(_03908_),
    .X(_03946_));
 sky130_fd_sc_hd__nand3_2 _11189_ (.A(_03771_),
    .B(_03754_),
    .C(_03756_),
    .Y(_03947_));
 sky130_fd_sc_hd__o21bai_1 _11190_ (.A1(_03781_),
    .A2(_03784_),
    .B1_N(_03782_),
    .Y(_03948_));
 sky130_fd_sc_hd__a22o_1 _11191_ (.A1(_00046_),
    .A2(_00530_),
    .B1(_06666_),
    .B2(_00049_),
    .X(_03949_));
 sky130_fd_sc_hd__nand4_1 _11192_ (.A(_00063_),
    .B(_00062_),
    .C(_05380_),
    .D(_05445_),
    .Y(_03950_));
 sky130_fd_sc_hd__a22o_1 _11193_ (.A1(_00058_),
    .A2(_05327_),
    .B1(_03949_),
    .B2(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__nand4_1 _11194_ (.A(_00444_),
    .B(_05327_),
    .C(_03949_),
    .D(_03950_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand3_1 _11195_ (.A(_03948_),
    .B(_03951_),
    .C(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__a21o_1 _11196_ (.A1(_03951_),
    .A2(_03952_),
    .B1(_03948_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(_03745_),
    .B(_03747_),
    .Y(_03955_));
 sky130_fd_sc_hd__a21o_1 _11198_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__nand3_1 _11199_ (.A(_03955_),
    .B(_03953_),
    .C(_03954_),
    .Y(_03957_));
 sky130_fd_sc_hd__a21bo_1 _11200_ (.A1(_03750_),
    .A2(_03749_),
    .B1_N(_03748_),
    .X(_03958_));
 sky130_fd_sc_hd__nand3_4 _11201_ (.A(_03956_),
    .B(_03957_),
    .C(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__a21o_1 _11202_ (.A1(_03956_),
    .A2(_03957_),
    .B1(_03958_),
    .X(_03961_));
 sky130_fd_sc_hd__a22oi_1 _11203_ (.A1(_00727_),
    .A2(_00197_),
    .B1(_00421_),
    .B2(_00728_),
    .Y(_03962_));
 sky130_fd_sc_hd__and4_1 _11204_ (.A(_01147_),
    .B(_01146_),
    .C(_04972_),
    .D(_05036_),
    .X(_03963_));
 sky130_fd_sc_hd__nor2_1 _11205_ (.A(_03962_),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand2_1 _11206_ (.A(_00077_),
    .B(_00550_),
    .Y(_03965_));
 sky130_fd_sc_hd__xnor2_1 _11207_ (.A(_03964_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__a22o_1 _11208_ (.A1(_00081_),
    .A2(_05187_),
    .B1(_05252_),
    .B2(_00086_),
    .X(_03967_));
 sky130_fd_sc_hd__nand4_1 _11209_ (.A(_00133_),
    .B(_03099_),
    .C(_05187_),
    .D(_05252_),
    .Y(_03968_));
 sky130_fd_sc_hd__and2_1 _11210_ (.A(_03152_),
    .B(_06623_),
    .X(_03969_));
 sky130_fd_sc_hd__nand3_1 _11211_ (.A(_03967_),
    .B(_03968_),
    .C(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hd__a21o_1 _11212_ (.A1(_03967_),
    .A2(_03968_),
    .B1(_03969_),
    .X(_03972_));
 sky130_fd_sc_hd__and2_2 _11213_ (.A(_00081_),
    .B(_05187_),
    .X(_03973_));
 sky130_fd_sc_hd__and2_2 _11214_ (.A(_00086_),
    .B(_06623_),
    .X(_03974_));
 sky130_fd_sc_hd__a32o_1 _11215_ (.A1(_03163_),
    .A2(_00421_),
    .A3(_03762_),
    .B1(_03973_),
    .B2(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__and3_1 _11216_ (.A(_03970_),
    .B(_03972_),
    .C(_03975_),
    .X(_03976_));
 sky130_fd_sc_hd__a21o_1 _11217_ (.A1(_03970_),
    .A2(_03972_),
    .B1(_03975_),
    .X(_03977_));
 sky130_fd_sc_hd__or2b_1 _11218_ (.A(_03976_),
    .B_N(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__xnor2_1 _11219_ (.A(_03966_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__a21oi_2 _11220_ (.A1(_03959_),
    .A2(_03961_),
    .B1(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__and3_1 _11221_ (.A(_03979_),
    .B(_03959_),
    .C(_03961_),
    .X(_03981_));
 sky130_fd_sc_hd__a211oi_4 _11222_ (.A1(_03796_),
    .A2(_03799_),
    .B1(_03980_),
    .C1(_03981_),
    .Y(_03983_));
 sky130_fd_sc_hd__o211a_1 _11223_ (.A1(_03980_),
    .A2(_03981_),
    .B1(_03796_),
    .C1(_03799_),
    .X(_03984_));
 sky130_fd_sc_hd__a211oi_4 _11224_ (.A1(_03754_),
    .A2(_03947_),
    .B1(_03983_),
    .C1(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__o211a_1 _11225_ (.A1(_03983_),
    .A2(_03984_),
    .B1(_03754_),
    .C1(_03947_),
    .X(_03986_));
 sky130_fd_sc_hd__nor4_1 _11226_ (.A(_03945_),
    .B(_03946_),
    .C(_03985_),
    .D(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__o22a_1 _11227_ (.A1(_03945_),
    .A2(_03946_),
    .B1(_03985_),
    .B2(_03986_),
    .X(_03988_));
 sky130_fd_sc_hd__a211o_2 _11228_ (.A1(_03812_),
    .A2(_03815_),
    .B1(_03987_),
    .C1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__o211ai_2 _11229_ (.A1(_03987_),
    .A2(_03988_),
    .B1(_03812_),
    .C1(_03815_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand4_4 _11230_ (.A(_03904_),
    .B(_03905_),
    .C(_03989_),
    .D(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__a22o_1 _11231_ (.A1(_03904_),
    .A2(_03905_),
    .B1(_03989_),
    .B2(_03990_),
    .X(_03992_));
 sky130_fd_sc_hd__o211a_1 _11232_ (.A1(_03816_),
    .A2(_03862_),
    .B1(_03991_),
    .C1(_03992_),
    .X(_03994_));
 sky130_fd_sc_hd__a211o_1 _11233_ (.A1(_03991_),
    .A2(_03992_),
    .B1(_03816_),
    .C1(_03862_),
    .X(_03995_));
 sky130_fd_sc_hd__and2b_1 _11234_ (.A_N(_03994_),
    .B(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__xnor2_4 _11235_ (.A(_03861_),
    .B(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__and2b_1 _11236_ (.A_N(_03822_),
    .B(_03819_),
    .X(_03998_));
 sky130_fd_sc_hd__a21oi_4 _11237_ (.A1(_03696_),
    .A2(_03823_),
    .B1(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__xnor2_4 _11238_ (.A(_03997_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__xnor2_1 _11239_ (.A(_03859_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__and2b_2 _11240_ (.A_N(_03827_),
    .B(_03824_),
    .X(_04002_));
 sky130_fd_sc_hd__a21oi_1 _11241_ (.A1(_03694_),
    .A2(_03828_),
    .B1(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_1 _11242_ (.A(_04001_),
    .B(_04003_),
    .Y(_04005_));
 sky130_fd_sc_hd__a21o_1 _11243_ (.A1(_03692_),
    .A2(_03693_),
    .B1(_03829_),
    .X(_04006_));
 sky130_fd_sc_hd__a31o_1 _11244_ (.A1(_03657_),
    .A2(_03667_),
    .A3(_04006_),
    .B1(_03832_),
    .X(_04007_));
 sky130_fd_sc_hd__or2_1 _11245_ (.A(_04005_),
    .B(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(_03133_),
    .B(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__a21oi_1 _11247_ (.A1(_04005_),
    .A2(_04007_),
    .B1(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__clkbuf_4 _11248_ (.A(_02707_),
    .X(_04011_));
 sky130_fd_sc_hd__o211a_1 _11249_ (.A1(_02129_),
    .A2(_01988_),
    .B1(_04011_),
    .C1(_02756_),
    .X(_04012_));
 sky130_fd_sc_hd__a221o_1 _11250_ (.A1(\MuI.result[6] ),
    .A2(_02739_),
    .B1(_02719_),
    .B2(_04391_),
    .C1(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__a32o_1 _11251_ (.A1(_02442_),
    .A2(_04327_),
    .A3(_02744_),
    .B1(_06045_),
    .B2(\FuI.Integer[6] ),
    .X(_04014_));
 sky130_fd_sc_hd__a2bb2o_1 _11252_ (.A1_N(_04327_),
    .A2_N(_02727_),
    .B1(_02945_),
    .B2(_04262_),
    .X(_04016_));
 sky130_fd_sc_hd__o21a_1 _11253_ (.A1(_02760_),
    .A2(_03838_),
    .B1(_02192_),
    .X(_04017_));
 sky130_fd_sc_hd__xor2_1 _11254_ (.A(_02757_),
    .B(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__a22o_1 _11255_ (.A1(\AuI.result[6] ),
    .A2(_02731_),
    .B1(_04018_),
    .B2(_02935_),
    .X(_04019_));
 sky130_fd_sc_hd__or3_1 _11256_ (.A(_04014_),
    .B(_04016_),
    .C(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__or2_1 _11257_ (.A(_04013_),
    .B(_04020_),
    .X(_04021_));
 sky130_fd_sc_hd__a311o_1 _11258_ (.A1(_02750_),
    .A2(_03855_),
    .A3(_03856_),
    .B1(_04010_),
    .C1(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__a31o_2 _11259_ (.A1(_02566_),
    .A2(_03315_),
    .A3(_03849_),
    .B1(_04022_),
    .X(net97));
 sky130_fd_sc_hd__or2_1 _11260_ (.A(_04001_),
    .B(_04003_),
    .X(_04023_));
 sky130_fd_sc_hd__nor2_1 _11261_ (.A(_03874_),
    .B(_03876_),
    .Y(_04024_));
 sky130_fd_sc_hd__a31o_1 _11262_ (.A1(_03820_),
    .A2(_04391_),
    .A3(_03877_),
    .B1(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__inv_2 _11263_ (.A(_03945_),
    .Y(_04026_));
 sky130_fd_sc_hd__or4_2 _11264_ (.A(_03945_),
    .B(_03946_),
    .C(_03985_),
    .D(_03986_),
    .X(_04027_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_03934_),
    .B(_03936_),
    .Y(_04028_));
 sky130_fd_sc_hd__a22oi_1 _11266_ (.A1(_00878_),
    .A2(_05649_),
    .B1(_03449_),
    .B2(_00877_),
    .Y(_04029_));
 sky130_fd_sc_hd__and4_1 _11267_ (.A(_00012_),
    .B(_00011_),
    .C(_03425_),
    .D(_05702_),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_1 _11268_ (.A(_04029_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_1 _11269_ (.A(_02840_),
    .B(_05585_),
    .Y(_04032_));
 sky130_fd_sc_hd__xnor2_1 _11270_ (.A(_04031_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a22oi_2 _11271_ (.A1(_02658_),
    .A2(_00783_),
    .B1(_05884_),
    .B2(_02593_),
    .Y(_04034_));
 sky130_fd_sc_hd__and4_1 _11272_ (.A(_06585_),
    .B(_06583_),
    .C(_00785_),
    .D(_00153_),
    .X(_04036_));
 sky130_fd_sc_hd__nand2_1 _11273_ (.A(_02712_),
    .B(_03247_),
    .Y(_04037_));
 sky130_fd_sc_hd__or3_1 _11274_ (.A(_04034_),
    .B(_04036_),
    .C(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__o21ai_1 _11275_ (.A1(_04034_),
    .A2(_04036_),
    .B1(_04037_),
    .Y(_04039_));
 sky130_fd_sc_hd__o21bai_1 _11276_ (.A1(_03927_),
    .A2(_03930_),
    .B1_N(_03929_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand3_1 _11277_ (.A(_04038_),
    .B(_04039_),
    .C(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__a21o_1 _11278_ (.A1(_04038_),
    .A2(_04039_),
    .B1(_04040_),
    .X(_04042_));
 sky130_fd_sc_hd__nand3_1 _11279_ (.A(_04033_),
    .B(_04041_),
    .C(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__a21o_1 _11280_ (.A1(_04041_),
    .A2(_04042_),
    .B1(_04033_),
    .X(_04044_));
 sky130_fd_sc_hd__nand3_2 _11281_ (.A(_03916_),
    .B(_04043_),
    .C(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__a21o_1 _11282_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_03916_),
    .X(_04047_));
 sky130_fd_sc_hd__nand3_2 _11283_ (.A(_04028_),
    .B(_04045_),
    .C(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__a21o_1 _11284_ (.A1(_04045_),
    .A2(_04047_),
    .B1(_04028_),
    .X(_04049_));
 sky130_fd_sc_hd__or4bb_2 _11285_ (.A(_03913_),
    .B(_03910_),
    .C_N(_04048_),
    .D_N(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__a2bb2o_1 _11286_ (.A1_N(_03913_),
    .A2_N(_03910_),
    .B1(_04048_),
    .B2(_04049_),
    .X(_04051_));
 sky130_fd_sc_hd__and3_1 _11287_ (.A(_03943_),
    .B(_04050_),
    .C(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__a21oi_1 _11288_ (.A1(_04050_),
    .A2(_04051_),
    .B1(_03943_),
    .Y(_04053_));
 sky130_fd_sc_hd__nand3_1 _11289_ (.A(_03979_),
    .B(_03959_),
    .C(_03961_),
    .Y(_04054_));
 sky130_fd_sc_hd__o21bai_1 _11290_ (.A1(_03922_),
    .A2(_03925_),
    .B1_N(_03923_),
    .Y(_04055_));
 sky130_fd_sc_hd__a22o_1 _11291_ (.A1(_00046_),
    .A2(_06666_),
    .B1(_00398_),
    .B2(_00049_),
    .X(_04056_));
 sky130_fd_sc_hd__nand4_1 _11292_ (.A(_00063_),
    .B(_00062_),
    .C(_05445_),
    .D(_05509_),
    .Y(_04058_));
 sky130_fd_sc_hd__a22o_1 _11293_ (.A1(_00058_),
    .A2(_05391_),
    .B1(_04056_),
    .B2(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__nand4_1 _11294_ (.A(_00444_),
    .B(_05391_),
    .C(_04056_),
    .D(_04058_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand3_1 _11295_ (.A(_04055_),
    .B(_04059_),
    .C(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a21o_1 _11296_ (.A1(_04059_),
    .A2(_04060_),
    .B1(_04055_),
    .X(_04062_));
 sky130_fd_sc_hd__nand2_1 _11297_ (.A(_03950_),
    .B(_03952_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21o_1 _11298_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__nand3_1 _11299_ (.A(_04063_),
    .B(_04061_),
    .C(_04062_),
    .Y(_04065_));
 sky130_fd_sc_hd__a21bo_1 _11300_ (.A1(_03955_),
    .A2(_03954_),
    .B1_N(_03953_),
    .X(_04066_));
 sky130_fd_sc_hd__nand3_2 _11301_ (.A(_04064_),
    .B(_04065_),
    .C(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a21o_1 _11302_ (.A1(_04064_),
    .A2(_04065_),
    .B1(_04066_),
    .X(_04069_));
 sky130_fd_sc_hd__a22oi_1 _11303_ (.A1(_00727_),
    .A2(_00421_),
    .B1(_00423_),
    .B2(_00728_),
    .Y(_04070_));
 sky130_fd_sc_hd__and4_1 _11304_ (.A(_03228_),
    .B(_03282_),
    .C(_05036_),
    .D(_00534_),
    .X(_04071_));
 sky130_fd_sc_hd__nor2_1 _11305_ (.A(_04070_),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _11306_ (.A(_00077_),
    .B(_00197_),
    .Y(_04073_));
 sky130_fd_sc_hd__xnor2_1 _11307_ (.A(_04072_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__a22oi_4 _11308_ (.A1(_00462_),
    .A2(_06518_),
    .B1(_06562_),
    .B2(_00086_),
    .Y(_04075_));
 sky130_fd_sc_hd__and4_2 _11309_ (.A(_00095_),
    .B(_00096_),
    .C(_05241_),
    .D(_05305_),
    .X(_04076_));
 sky130_fd_sc_hd__nand2_1 _11310_ (.A(_00088_),
    .B(_05187_),
    .Y(_04077_));
 sky130_fd_sc_hd__or3_1 _11311_ (.A(_04075_),
    .B(_04076_),
    .C(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__o21ai_1 _11312_ (.A1(_04075_),
    .A2(_04076_),
    .B1(_04077_),
    .Y(_04080_));
 sky130_fd_sc_hd__a21bo_1 _11313_ (.A1(_03967_),
    .A2(_03969_),
    .B1_N(_03968_),
    .X(_04081_));
 sky130_fd_sc_hd__and3_1 _11314_ (.A(_04078_),
    .B(_04080_),
    .C(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__a21o_1 _11315_ (.A1(_04078_),
    .A2(_04080_),
    .B1(_04081_),
    .X(_04083_));
 sky130_fd_sc_hd__and2b_1 _11316_ (.A_N(_04082_),
    .B(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__xor2_1 _11317_ (.A(_04074_),
    .B(_04084_),
    .X(_04085_));
 sky130_fd_sc_hd__a21oi_2 _11318_ (.A1(_04067_),
    .A2(_04069_),
    .B1(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__and3_1 _11319_ (.A(_04085_),
    .B(_04067_),
    .C(_04069_),
    .X(_04087_));
 sky130_fd_sc_hd__a211oi_4 _11320_ (.A1(_03938_),
    .A2(_03941_),
    .B1(_04086_),
    .C1(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__o211a_1 _11321_ (.A1(_04086_),
    .A2(_04087_),
    .B1(_03938_),
    .C1(_03941_),
    .X(_04089_));
 sky130_fd_sc_hd__a211oi_4 _11322_ (.A1(_03959_),
    .A2(_04054_),
    .B1(_04088_),
    .C1(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__o211a_1 _11323_ (.A1(_04088_),
    .A2(_04089_),
    .B1(_03959_),
    .C1(_04054_),
    .X(_04091_));
 sky130_fd_sc_hd__o22a_1 _11324_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04090_),
    .B2(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__nor4_2 _11325_ (.A(_04052_),
    .B(_04053_),
    .C(_04090_),
    .D(_04091_),
    .Y(_04093_));
 sky130_fd_sc_hd__a211o_2 _11326_ (.A1(_04026_),
    .A2(_04027_),
    .B1(_04092_),
    .C1(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__o211ai_4 _11327_ (.A1(_04092_),
    .A2(_04093_),
    .B1(_04026_),
    .C1(_04027_),
    .Y(_04095_));
 sky130_fd_sc_hd__inv_2 _11328_ (.A(_03898_),
    .Y(_04096_));
 sky130_fd_sc_hd__and3_1 _11329_ (.A(_03879_),
    .B(_03898_),
    .C(_03899_),
    .X(_04097_));
 sky130_fd_sc_hd__and3_1 _11330_ (.A(_00506_),
    .B(_00676_),
    .C(_00048_),
    .X(_04098_));
 sky130_fd_sc_hd__a22o_1 _11331_ (.A1(_00676_),
    .A2(_00048_),
    .B1(_00040_),
    .B2(_00506_),
    .X(_04099_));
 sky130_fd_sc_hd__a21bo_1 _11332_ (.A1(_04725_),
    .A2(_04098_),
    .B1_N(_04099_),
    .X(_04101_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(_02965_),
    .B(_04596_),
    .Y(_04102_));
 sky130_fd_sc_hd__xor2_4 _11334_ (.A(_04101_),
    .B(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__a32o_2 _11335_ (.A1(_03525_),
    .A2(_04531_),
    .A3(_03866_),
    .B1(_03865_),
    .B2(_04660_),
    .X(_04104_));
 sky130_fd_sc_hd__xor2_4 _11336_ (.A(_04103_),
    .B(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__and2_2 _11337_ (.A(_06429_),
    .B(_04531_),
    .X(_04106_));
 sky130_fd_sc_hd__xnor2_4 _11338_ (.A(_04105_),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__and2_1 _11339_ (.A(_03869_),
    .B(_03870_),
    .X(_04108_));
 sky130_fd_sc_hd__a21oi_2 _11340_ (.A1(_03871_),
    .A2(_03872_),
    .B1(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__xor2_4 _11341_ (.A(_04107_),
    .B(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__nand2_1 _11342_ (.A(_00502_),
    .B(_04467_),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_4 _11343_ (.A(_04110_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a211oi_2 _11344_ (.A1(_03721_),
    .A2(_03726_),
    .B1(_03893_),
    .C1(_03894_),
    .Y(_04114_));
 sky130_fd_sc_hd__a21o_1 _11345_ (.A1(_03966_),
    .A2(_03977_),
    .B1(_03976_),
    .X(_04115_));
 sky130_fd_sc_hd__o21bai_1 _11346_ (.A1(_03962_),
    .A2(_03965_),
    .B1_N(_03963_),
    .Y(_04116_));
 sky130_fd_sc_hd__a22o_1 _11347_ (.A1(_02980_),
    .A2(_00445_),
    .B1(_04907_),
    .B2(_02983_),
    .X(_04117_));
 sky130_fd_sc_hd__nand4_1 _11348_ (.A(_03389_),
    .B(_02984_),
    .C(_00445_),
    .D(_00550_),
    .Y(_04118_));
 sky130_fd_sc_hd__a22o_1 _11349_ (.A1(_00345_),
    .A2(_06613_),
    .B1(_04117_),
    .B2(_04118_),
    .X(_04119_));
 sky130_fd_sc_hd__nand4_1 _11350_ (.A(_02987_),
    .B(_06613_),
    .C(_04117_),
    .D(_04118_),
    .Y(_04120_));
 sky130_fd_sc_hd__nand3_2 _11351_ (.A(_04116_),
    .B(_04119_),
    .C(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__a21o_1 _11352_ (.A1(_04119_),
    .A2(_04120_),
    .B1(_04116_),
    .X(_04123_));
 sky130_fd_sc_hd__nand2_1 _11353_ (.A(_03885_),
    .B(_03887_),
    .Y(_04124_));
 sky130_fd_sc_hd__a21o_1 _11354_ (.A1(_04121_),
    .A2(_04123_),
    .B1(_04124_),
    .X(_04125_));
 sky130_fd_sc_hd__nand3_2 _11355_ (.A(_04124_),
    .B(_04121_),
    .C(_04123_),
    .Y(_04126_));
 sky130_fd_sc_hd__and3_1 _11356_ (.A(_04115_),
    .B(_04125_),
    .C(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__a21oi_1 _11357_ (.A1(_04125_),
    .A2(_04126_),
    .B1(_04115_),
    .Y(_04128_));
 sky130_fd_sc_hd__a211o_1 _11358_ (.A1(_03888_),
    .A2(_03892_),
    .B1(_04127_),
    .C1(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__o211ai_1 _11359_ (.A1(_04127_),
    .A2(_04128_),
    .B1(_03888_),
    .C1(_03892_),
    .Y(_04130_));
 sky130_fd_sc_hd__o211ai_2 _11360_ (.A1(_03893_),
    .A2(_04114_),
    .B1(_04129_),
    .C1(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__a211o_1 _11361_ (.A1(_04129_),
    .A2(_04130_),
    .B1(_03893_),
    .C1(_04114_),
    .X(_04132_));
 sky130_fd_sc_hd__nand3_1 _11362_ (.A(_04113_),
    .B(_04131_),
    .C(_04132_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21o_1 _11363_ (.A1(_04131_),
    .A2(_04132_),
    .B1(_04113_),
    .X(_04135_));
 sky130_fd_sc_hd__o211ai_4 _11364_ (.A1(_03983_),
    .A2(_03985_),
    .B1(_04134_),
    .C1(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__a211o_1 _11365_ (.A1(_04134_),
    .A2(_04135_),
    .B1(_03983_),
    .C1(_03985_),
    .X(_04137_));
 sky130_fd_sc_hd__o211ai_4 _11366_ (.A1(_04096_),
    .A2(_04097_),
    .B1(_04136_),
    .C1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a211o_1 _11367_ (.A1(_04136_),
    .A2(_04137_),
    .B1(_04096_),
    .C1(_04097_),
    .X(_04139_));
 sky130_fd_sc_hd__and4_1 _11368_ (.A(_04094_),
    .B(_04095_),
    .C(_04138_),
    .D(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__a22oi_4 _11369_ (.A1(_04094_),
    .A2(_04095_),
    .B1(_04138_),
    .B2(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__a211oi_4 _11370_ (.A1(_03989_),
    .A2(_03991_),
    .B1(_04140_),
    .C1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__o211a_1 _11371_ (.A1(_04140_),
    .A2(_04141_),
    .B1(_03989_),
    .C1(_03991_),
    .X(_04143_));
 sky130_fd_sc_hd__a211oi_4 _11372_ (.A1(_03902_),
    .A2(_03904_),
    .B1(_04142_),
    .C1(_04143_),
    .Y(_04145_));
 sky130_fd_sc_hd__o211a_1 _11373_ (.A1(_04142_),
    .A2(_04143_),
    .B1(_03902_),
    .C1(_03904_),
    .X(_04146_));
 sky130_fd_sc_hd__nor2_2 _11374_ (.A(_04145_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__a21oi_2 _11375_ (.A1(_03861_),
    .A2(_03995_),
    .B1(_03994_),
    .Y(_04148_));
 sky130_fd_sc_hd__xnor2_4 _11376_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__xnor2_1 _11377_ (.A(_04025_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__nor2_2 _11378_ (.A(_03997_),
    .B(_03999_),
    .Y(_04151_));
 sky130_fd_sc_hd__o21ba_1 _11379_ (.A1(_03859_),
    .A2(_04000_),
    .B1_N(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__xnor2_1 _11380_ (.A(_04150_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__a21oi_1 _11381_ (.A1(_04023_),
    .A2(_04008_),
    .B1(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__and3_1 _11382_ (.A(_04023_),
    .B(_04008_),
    .C(_04153_),
    .X(_04155_));
 sky130_fd_sc_hd__or2_1 _11383_ (.A(_04154_),
    .B(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__or2_1 _11384_ (.A(_02566_),
    .B(_02568_),
    .X(_04157_));
 sky130_fd_sc_hd__or3b_1 _11385_ (.A(_02709_),
    .B(_02064_),
    .C_N(_06023_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_4 _11386_ (.A(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__a21oi_1 _11387_ (.A1(_02566_),
    .A2(_02568_),
    .B1(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__buf_4 _11388_ (.A(_02935_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _11389_ (.A(_02771_),
    .B(_02772_),
    .Y(_04162_));
 sky130_fd_sc_hd__o21a_1 _11390_ (.A1(_02757_),
    .A2(_04017_),
    .B1(_01988_),
    .X(_04163_));
 sky130_fd_sc_hd__xnor2_1 _11391_ (.A(_04162_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__a2bb2o_1 _11392_ (.A1_N(_04391_),
    .A2_N(_02728_),
    .B1(_04162_),
    .B2(_03494_),
    .X(_04166_));
 sky130_fd_sc_hd__o21a_1 _11393_ (.A1(_02496_),
    .A2(_04391_),
    .B1(_02722_),
    .X(_04167_));
 sky130_fd_sc_hd__and3_1 _11394_ (.A(_02496_),
    .B(_04391_),
    .C(_02743_),
    .X(_04168_));
 sky130_fd_sc_hd__a221o_1 _11395_ (.A1(\MuI.result[7] ),
    .A2(_02737_),
    .B1(_02945_),
    .B2(_04327_),
    .C1(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__a221o_1 _11396_ (.A1(_04467_),
    .A2(_03675_),
    .B1(_02938_),
    .B2(\AuI.result[7] ),
    .C1(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__a2111o_1 _11397_ (.A1(\FuI.Integer[7] ),
    .A2(_06056_),
    .B1(_04166_),
    .C1(_04167_),
    .D1(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__a21o_1 _11398_ (.A1(_04161_),
    .A2(_04164_),
    .B1(_04171_),
    .X(_04172_));
 sky130_fd_sc_hd__a21oi_2 _11399_ (.A1(_04157_),
    .A2(_04160_),
    .B1(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__or2b_1 _11400_ (.A(_04327_),
    .B_N(_02442_),
    .X(_04174_));
 sky130_fd_sc_hd__o31ai_1 _11401_ (.A1(_02887_),
    .A2(_02759_),
    .A3(_03850_),
    .B1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__a31o_1 _11402_ (.A1(_02879_),
    .A2(_02886_),
    .A3(_02757_),
    .B1(_02887_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(_04175_),
    .A1(_04177_),
    .S(_02926_),
    .X(_04178_));
 sky130_fd_sc_hd__o21ai_1 _11404_ (.A1(_02773_),
    .A2(_04178_),
    .B1(_02750_),
    .Y(_04179_));
 sky130_fd_sc_hd__a21o_1 _11405_ (.A1(_02773_),
    .A2(_04178_),
    .B1(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__o211ai_4 _11406_ (.A1(_06428_),
    .A2(_04156_),
    .B1(_04173_),
    .C1(_04180_),
    .Y(net98));
 sky130_fd_sc_hd__and3_1 _11407_ (.A(_03809_),
    .B(_04467_),
    .C(_04110_),
    .X(_04181_));
 sky130_fd_sc_hd__o21ba_1 _11408_ (.A1(_04107_),
    .A2(_04109_),
    .B1_N(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__nand4_2 _11409_ (.A(_04094_),
    .B(_04095_),
    .C(_04138_),
    .D(_04139_),
    .Y(_04183_));
 sky130_fd_sc_hd__inv_2 _11410_ (.A(_04052_),
    .Y(_04184_));
 sky130_fd_sc_hd__or4_2 _11411_ (.A(_04052_),
    .B(_04053_),
    .C(_04090_),
    .D(_04091_),
    .X(_04185_));
 sky130_fd_sc_hd__nand3_1 _11412_ (.A(_04085_),
    .B(_04067_),
    .C(_04069_),
    .Y(_04187_));
 sky130_fd_sc_hd__o21bai_1 _11413_ (.A1(_04029_),
    .A2(_04032_),
    .B1_N(_04030_),
    .Y(_04188_));
 sky130_fd_sc_hd__a22o_1 _11414_ (.A1(_00216_),
    .A2(_03051_),
    .B1(_05574_),
    .B2(_00217_),
    .X(_04189_));
 sky130_fd_sc_hd__nand4_1 _11415_ (.A(_02905_),
    .B(_02959_),
    .C(_03051_),
    .D(_03071_),
    .Y(_04190_));
 sky130_fd_sc_hd__a22o_1 _11416_ (.A1(_00221_),
    .A2(_05456_),
    .B1(_04189_),
    .B2(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__nand4_1 _11417_ (.A(_03013_),
    .B(_05456_),
    .C(_04189_),
    .D(_04190_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand3_1 _11418_ (.A(_04188_),
    .B(_04191_),
    .C(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__a21o_1 _11419_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_04188_),
    .X(_04194_));
 sky130_fd_sc_hd__nand2_1 _11420_ (.A(_04058_),
    .B(_04060_),
    .Y(_04195_));
 sky130_fd_sc_hd__a21o_1 _11421_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__nand3_1 _11422_ (.A(_04195_),
    .B(_04193_),
    .C(_04194_),
    .Y(_04198_));
 sky130_fd_sc_hd__a21bo_1 _11423_ (.A1(_04063_),
    .A2(_04062_),
    .B1_N(_04061_),
    .X(_04199_));
 sky130_fd_sc_hd__nand3_2 _11424_ (.A(_04196_),
    .B(_04198_),
    .C(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__a21o_1 _11425_ (.A1(_04196_),
    .A2(_04198_),
    .B1(_04199_),
    .X(_04201_));
 sky130_fd_sc_hd__a22oi_1 _11426_ (.A1(_00727_),
    .A2(_00423_),
    .B1(_05198_),
    .B2(_00728_),
    .Y(_04202_));
 sky130_fd_sc_hd__and4_1 _11427_ (.A(_03228_),
    .B(_03282_),
    .C(_00534_),
    .D(_06525_),
    .X(_04203_));
 sky130_fd_sc_hd__nor2_1 _11428_ (.A(_04202_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_1 _11429_ (.A(_03324_),
    .B(_05047_),
    .Y(_04205_));
 sky130_fd_sc_hd__xnor2_1 _11430_ (.A(_04204_),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nor3_1 _11431_ (.A(_04075_),
    .B(_04076_),
    .C(_04077_),
    .Y(_04207_));
 sky130_fd_sc_hd__a22oi_1 _11432_ (.A1(_00132_),
    .A2(_05316_),
    .B1(_05380_),
    .B2(_00133_),
    .Y(_04209_));
 sky130_fd_sc_hd__and4_1 _11433_ (.A(_00086_),
    .B(_00081_),
    .C(_00412_),
    .D(_00530_),
    .X(_04210_));
 sky130_fd_sc_hd__nand2_4 _11434_ (.A(_00088_),
    .B(_06568_),
    .Y(_04211_));
 sky130_fd_sc_hd__o21ai_1 _11435_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__or3_1 _11436_ (.A(_04211_),
    .B(_04209_),
    .C(_04210_),
    .X(_04213_));
 sky130_fd_sc_hd__o211a_1 _11437_ (.A1(_04076_),
    .A2(_04207_),
    .B1(_04212_),
    .C1(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__a211o_1 _11438_ (.A1(_04212_),
    .A2(_04213_),
    .B1(_04076_),
    .C1(_04207_),
    .X(_04215_));
 sky130_fd_sc_hd__or2b_1 _11439_ (.A(_04214_),
    .B_N(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__xnor2_1 _11440_ (.A(_04206_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__a21oi_1 _11441_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__and3_1 _11442_ (.A(_04217_),
    .B(_04200_),
    .C(_04201_),
    .X(_04219_));
 sky130_fd_sc_hd__a211oi_1 _11443_ (.A1(_04045_),
    .A2(_04048_),
    .B1(_04218_),
    .C1(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__o211a_1 _11444_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04045_),
    .C1(_04048_),
    .X(_04221_));
 sky130_fd_sc_hd__a211o_1 _11445_ (.A1(_04067_),
    .A2(_04187_),
    .B1(_04220_),
    .C1(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__o211ai_2 _11446_ (.A1(_04220_),
    .A2(_04221_),
    .B1(_04067_),
    .C1(_04187_),
    .Y(_04223_));
 sky130_fd_sc_hd__a22o_1 _11447_ (.A1(_02658_),
    .A2(_03082_),
    .B1(_00789_),
    .B2(_06585_),
    .X(_04224_));
 sky130_fd_sc_hd__nand4_2 _11448_ (.A(_02593_),
    .B(_02658_),
    .C(_03082_),
    .D(_00789_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand4_1 _11449_ (.A(_06620_),
    .B(_03257_),
    .C(_04224_),
    .D(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__a22o_1 _11450_ (.A1(_06620_),
    .A2(_03257_),
    .B1(_04224_),
    .B2(_04225_),
    .X(_04227_));
 sky130_fd_sc_hd__o21bai_1 _11451_ (.A1(_04034_),
    .A2(_04037_),
    .B1_N(_04036_),
    .Y(_04228_));
 sky130_fd_sc_hd__and3_1 _11452_ (.A(_04226_),
    .B(_04227_),
    .C(_04228_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_1 _11453_ (.A1(_04226_),
    .A2(_04227_),
    .B1(_04228_),
    .Y(_04231_));
 sky130_fd_sc_hd__a22oi_1 _11454_ (.A1(_00878_),
    .A2(_05702_),
    .B1(_05767_),
    .B2(_00877_),
    .Y(_04232_));
 sky130_fd_sc_hd__and4_1 _11455_ (.A(_06606_),
    .B(_06601_),
    .C(_06537_),
    .D(_00385_),
    .X(_04233_));
 sky130_fd_sc_hd__nor2_1 _11456_ (.A(_04232_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _11457_ (.A(_02840_),
    .B(_05649_),
    .Y(_04235_));
 sky130_fd_sc_hd__xnor2_1 _11458_ (.A(_04234_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__or3b_1 _11459_ (.A(_04230_),
    .B(_04231_),
    .C_N(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__o21bai_1 _11460_ (.A1(_04230_),
    .A2(_04231_),
    .B1_N(_04236_),
    .Y(_04238_));
 sky130_fd_sc_hd__nor2_1 _11461_ (.A(_03909_),
    .B(_03910_),
    .Y(_04239_));
 sky130_fd_sc_hd__a21o_1 _11462_ (.A1(_04237_),
    .A2(_04238_),
    .B1(_04239_),
    .X(_04241_));
 sky130_fd_sc_hd__nand3_1 _11463_ (.A(_04239_),
    .B(_04237_),
    .C(_04238_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2_1 _11464_ (.A(_04041_),
    .B(_04043_),
    .Y(_04243_));
 sky130_fd_sc_hd__and3_1 _11465_ (.A(_04241_),
    .B(_04242_),
    .C(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__a21oi_1 _11466_ (.A1(_04241_),
    .A2(_04242_),
    .B1(_04243_),
    .Y(_04245_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(_04244_),
    .B(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__xor2_1 _11468_ (.A(_04050_),
    .B(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__a21oi_2 _11469_ (.A1(_04222_),
    .A2(_04223_),
    .B1(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__and3_2 _11470_ (.A(_04247_),
    .B(_04222_),
    .C(_04223_),
    .X(_04249_));
 sky130_fd_sc_hd__a211o_2 _11471_ (.A1(_04184_),
    .A2(_04185_),
    .B1(_04248_),
    .C1(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__o211ai_4 _11472_ (.A1(_04248_),
    .A2(_04249_),
    .B1(_04184_),
    .C1(_04185_),
    .Y(_04252_));
 sky130_fd_sc_hd__inv_2 _11473_ (.A(_04131_),
    .Y(_04253_));
 sky130_fd_sc_hd__and3_1 _11474_ (.A(_04113_),
    .B(_04131_),
    .C(_04132_),
    .X(_04254_));
 sky130_fd_sc_hd__and3_1 _11475_ (.A(_06434_),
    .B(_03604_),
    .C(_00033_),
    .X(_04255_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(_03604_),
    .A2(_00033_),
    .B1(_06612_),
    .B2(_06434_),
    .X(_04256_));
 sky130_fd_sc_hd__a21bo_1 _11477_ (.A1(_06613_),
    .A2(_04255_),
    .B1_N(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_1 _11478_ (.A(_02965_),
    .B(_04660_),
    .Y(_04258_));
 sky130_fd_sc_hd__xor2_2 _11479_ (.A(_04257_),
    .B(_04258_),
    .X(_04259_));
 sky130_fd_sc_hd__a32o_1 _11480_ (.A1(_03525_),
    .A2(_04596_),
    .A3(_04099_),
    .B1(_04098_),
    .B2(_04725_),
    .X(_04260_));
 sky130_fd_sc_hd__xor2_2 _11481_ (.A(_04259_),
    .B(_04260_),
    .X(_04261_));
 sky130_fd_sc_hd__and2_1 _11482_ (.A(_03722_),
    .B(_04596_),
    .X(_04263_));
 sky130_fd_sc_hd__xnor2_2 _11483_ (.A(_04261_),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__and2_1 _11484_ (.A(_04103_),
    .B(_04104_),
    .X(_04265_));
 sky130_fd_sc_hd__a21oi_2 _11485_ (.A1(_04105_),
    .A2(_04106_),
    .B1(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__xor2_4 _11486_ (.A(_04264_),
    .B(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__nand2_1 _11487_ (.A(_00502_),
    .B(_04542_),
    .Y(_04268_));
 sky130_fd_sc_hd__xnor2_4 _11488_ (.A(_04267_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__a211oi_1 _11489_ (.A1(_03888_),
    .A2(_03892_),
    .B1(_04127_),
    .C1(_04128_),
    .Y(_04270_));
 sky130_fd_sc_hd__a21o_1 _11490_ (.A1(_04074_),
    .A2(_04083_),
    .B1(_04082_),
    .X(_04271_));
 sky130_fd_sc_hd__o21bai_1 _11491_ (.A1(_04070_),
    .A2(_04073_),
    .B1_N(_04071_),
    .Y(_04272_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(_02980_),
    .A2(_04907_),
    .B1(_04972_),
    .B2(_00281_),
    .X(_04274_));
 sky130_fd_sc_hd__nand4_1 _11493_ (.A(_02983_),
    .B(_02984_),
    .C(_00550_),
    .D(_04972_),
    .Y(_04275_));
 sky130_fd_sc_hd__a22o_1 _11494_ (.A1(_00345_),
    .A2(_04854_),
    .B1(_04274_),
    .B2(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__nand4_1 _11495_ (.A(_02987_),
    .B(_04854_),
    .C(_04274_),
    .D(_04275_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand3_2 _11496_ (.A(_04272_),
    .B(_04276_),
    .C(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__a21o_1 _11497_ (.A1(_04276_),
    .A2(_04277_),
    .B1(_04272_),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_1 _11498_ (.A(_04118_),
    .B(_04120_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21o_1 _11499_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__nand3_2 _11500_ (.A(_04280_),
    .B(_04278_),
    .C(_04279_),
    .Y(_04282_));
 sky130_fd_sc_hd__and3_1 _11501_ (.A(_04271_),
    .B(_04281_),
    .C(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__a21oi_1 _11502_ (.A1(_04281_),
    .A2(_04282_),
    .B1(_04271_),
    .Y(_04284_));
 sky130_fd_sc_hd__a211o_1 _11503_ (.A1(_04121_),
    .A2(_04126_),
    .B1(_04283_),
    .C1(_04284_),
    .X(_04285_));
 sky130_fd_sc_hd__o211ai_1 _11504_ (.A1(_04283_),
    .A2(_04284_),
    .B1(_04121_),
    .C1(_04126_),
    .Y(_04286_));
 sky130_fd_sc_hd__o211ai_2 _11505_ (.A1(_04127_),
    .A2(_04270_),
    .B1(_04285_),
    .C1(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__a211o_1 _11506_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04127_),
    .C1(_04270_),
    .X(_04288_));
 sky130_fd_sc_hd__nand3_1 _11507_ (.A(_04269_),
    .B(_04287_),
    .C(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__a21o_1 _11508_ (.A1(_04287_),
    .A2(_04288_),
    .B1(_04269_),
    .X(_04290_));
 sky130_fd_sc_hd__o211ai_4 _11509_ (.A1(_04088_),
    .A2(_04090_),
    .B1(_04289_),
    .C1(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a211o_1 _11510_ (.A1(_04289_),
    .A2(_04290_),
    .B1(_04088_),
    .C1(_04090_),
    .X(_04292_));
 sky130_fd_sc_hd__o211ai_4 _11511_ (.A1(_04253_),
    .A2(_04254_),
    .B1(_04291_),
    .C1(_04292_),
    .Y(_04293_));
 sky130_fd_sc_hd__a211o_1 _11512_ (.A1(_04291_),
    .A2(_04292_),
    .B1(_04253_),
    .C1(_04254_),
    .X(_04295_));
 sky130_fd_sc_hd__and4_1 _11513_ (.A(_04250_),
    .B(_04252_),
    .C(_04293_),
    .D(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__a22oi_4 _11514_ (.A1(_04250_),
    .A2(_04252_),
    .B1(_04293_),
    .B2(_04295_),
    .Y(_04297_));
 sky130_fd_sc_hd__a211oi_4 _11515_ (.A1(_04094_),
    .A2(_04183_),
    .B1(_04296_),
    .C1(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_1 _11516_ (.A1(_04296_),
    .A2(_04297_),
    .B1(_04094_),
    .C1(_04183_),
    .X(_04299_));
 sky130_fd_sc_hd__a211o_1 _11517_ (.A1(_04136_),
    .A2(_04138_),
    .B1(_04298_),
    .C1(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__o211ai_2 _11518_ (.A1(_04298_),
    .A2(_04299_),
    .B1(_04136_),
    .C1(_04138_),
    .Y(_04301_));
 sky130_fd_sc_hd__o211a_2 _11519_ (.A1(_04142_),
    .A2(_04145_),
    .B1(_04300_),
    .C1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__a211oi_4 _11520_ (.A1(_04300_),
    .A2(_04301_),
    .B1(_04142_),
    .C1(_04145_),
    .Y(_04303_));
 sky130_fd_sc_hd__or3_1 _11521_ (.A(_04182_),
    .B(_04302_),
    .C(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__o21ai_1 _11522_ (.A1(_04302_),
    .A2(_04303_),
    .B1(_04182_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand2_1 _11523_ (.A(_04304_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__and2b_2 _11524_ (.A_N(_04148_),
    .B(_04147_),
    .X(_04308_));
 sky130_fd_sc_hd__a21oi_1 _11525_ (.A1(_04025_),
    .A2(_04149_),
    .B1(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__or2_1 _11526_ (.A(_04307_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__nand2_1 _11527_ (.A(_04307_),
    .B(_04309_),
    .Y(_04311_));
 sky130_fd_sc_hd__and2_1 _11528_ (.A(_04310_),
    .B(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__nor2_1 _11529_ (.A(_04005_),
    .B(_04153_),
    .Y(_04313_));
 sky130_fd_sc_hd__and3b_1 _11530_ (.A_N(_03660_),
    .B(_03833_),
    .C(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__and3_1 _11531_ (.A(_03295_),
    .B(_03661_),
    .C(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__and2_1 _11532_ (.A(_04150_),
    .B(_04152_),
    .X(_04317_));
 sky130_fd_sc_hd__o21a_1 _11533_ (.A1(_04150_),
    .A2(_04152_),
    .B1(_04023_),
    .X(_04318_));
 sky130_fd_sc_hd__a21oi_1 _11534_ (.A1(_03657_),
    .A2(_04006_),
    .B1(_03832_),
    .Y(_04319_));
 sky130_fd_sc_hd__a2bb2o_1 _11535_ (.A1_N(_04317_),
    .A2_N(_04318_),
    .B1(_04313_),
    .B2(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__a21o_1 _11536_ (.A1(_03664_),
    .A2(_04314_),
    .B1(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__a21oi_2 _11537_ (.A1(_02703_),
    .A2(_04315_),
    .B1(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__or2b_1 _11538_ (.A(_04312_),
    .B_N(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__or2b_1 _11539_ (.A(_04322_),
    .B_N(_04312_),
    .X(_04324_));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(_02786_),
    .Y(_04325_));
 sky130_fd_sc_hd__o21a_1 _11541_ (.A1(_02773_),
    .A2(_04163_),
    .B1(_01891_),
    .X(_04326_));
 sky130_fd_sc_hd__xnor2_1 _11542_ (.A(_04325_),
    .B(_04326_),
    .Y(_04328_));
 sky130_fd_sc_hd__a2bb2o_1 _11543_ (.A1_N(_04467_),
    .A2_N(_02728_),
    .B1(_02938_),
    .B2(\AuI.result[8] ),
    .X(_04329_));
 sky130_fd_sc_hd__a32o_1 _11544_ (.A1(_02550_),
    .A2(_04467_),
    .A3(_02743_),
    .B1(_02944_),
    .B2(_04391_),
    .X(_04330_));
 sky130_fd_sc_hd__a221o_1 _11545_ (.A1(\MuI.result[8] ),
    .A2(_02737_),
    .B1(_04011_),
    .B2(_04325_),
    .C1(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__a221o_1 _11546_ (.A1(\FuI.Integer[8] ),
    .A2(_02931_),
    .B1(_02719_),
    .B2(_04542_),
    .C1(_04331_),
    .X(_04332_));
 sky130_fd_sc_hd__a211o_1 _11547_ (.A1(_02550_),
    .A2(_02724_),
    .B1(_04329_),
    .C1(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__a21bo_1 _11548_ (.A1(_02546_),
    .A2(_02569_),
    .B1_N(_04157_),
    .X(_04334_));
 sky130_fd_sc_hd__and3b_1 _11549_ (.A_N(_02570_),
    .B(_02741_),
    .C(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__a211o_1 _11550_ (.A1(_04161_),
    .A2(_04328_),
    .B1(_04333_),
    .C1(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(_02772_),
    .B(_02889_),
    .Y(_04337_));
 sky130_fd_sc_hd__xnor2_1 _11552_ (.A(_04325_),
    .B(_04337_),
    .Y(_04339_));
 sky130_fd_sc_hd__or2b_1 _11553_ (.A(_02924_),
    .B_N(_02775_),
    .X(_04340_));
 sky130_fd_sc_hd__a21oi_1 _11554_ (.A1(_04339_),
    .A2(_04340_),
    .B1(_02713_),
    .Y(_04341_));
 sky130_fd_sc_hd__o21a_1 _11555_ (.A1(_04339_),
    .A2(_04340_),
    .B1(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__a311o_2 _11556_ (.A1(_03134_),
    .A2(_04323_),
    .A3(_04324_),
    .B1(_04336_),
    .C1(_04342_),
    .X(net99));
 sky130_fd_sc_hd__a21boi_1 _11557_ (.A1(_02771_),
    .A2(_04175_),
    .B1_N(_02772_),
    .Y(_04343_));
 sky130_fd_sc_hd__o21bai_1 _11558_ (.A1(_02784_),
    .A2(_04343_),
    .B1_N(_02785_),
    .Y(_04344_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(_04344_),
    .A1(_02890_),
    .S(_02928_),
    .X(_04345_));
 sky130_fd_sc_hd__xnor2_2 _11560_ (.A(_02790_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__xnor2_1 _11561_ (.A(_02546_),
    .B(_02548_),
    .Y(_04347_));
 sky130_fd_sc_hd__nor2_1 _11562_ (.A(_02570_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__o21a_1 _11563_ (.A1(_02786_),
    .A2(_04326_),
    .B1(_01702_),
    .X(_04349_));
 sky130_fd_sc_hd__xor2_1 _11564_ (.A(_02790_),
    .B(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__a2bb2o_1 _11565_ (.A1_N(_04542_),
    .A2_N(_02728_),
    .B1(_02938_),
    .B2(\AuI.result[9] ),
    .X(_04351_));
 sky130_fd_sc_hd__a32o_1 _11566_ (.A1(_02604_),
    .A2(_04542_),
    .A3(_02744_),
    .B1(_02945_),
    .B2(_04467_),
    .X(_04352_));
 sky130_fd_sc_hd__a2bb2o_1 _11567_ (.A1_N(_03306_),
    .A2_N(_02790_),
    .B1(\MuI.result[9] ),
    .B2(_02737_),
    .X(_04353_));
 sky130_fd_sc_hd__a22o_1 _11568_ (.A1(\FuI.Integer[9] ),
    .A2(_06045_),
    .B1(_02718_),
    .B2(_04607_),
    .X(_04354_));
 sky130_fd_sc_hd__or3_1 _11569_ (.A(_04352_),
    .B(_04353_),
    .C(_04354_),
    .X(_04355_));
 sky130_fd_sc_hd__a211o_1 _11570_ (.A1(_02604_),
    .A2(_02724_),
    .B1(_04351_),
    .C1(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_1 _11571_ (.A1(_04161_),
    .A2(_04350_),
    .B1(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_04310_),
    .B(_04324_),
    .Y(_04359_));
 sky130_fd_sc_hd__inv_2 _11573_ (.A(_04302_),
    .Y(_04360_));
 sky130_fd_sc_hd__or2_1 _11574_ (.A(_04264_),
    .B(_04266_),
    .X(_04361_));
 sky130_fd_sc_hd__nand3_1 _11575_ (.A(_03831_),
    .B(_04542_),
    .C(_04267_),
    .Y(_04362_));
 sky130_fd_sc_hd__a211oi_2 _11576_ (.A1(_04136_),
    .A2(_04138_),
    .B1(_04298_),
    .C1(_04299_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand4_2 _11577_ (.A(_04250_),
    .B(_04252_),
    .C(_04293_),
    .D(_04295_),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_1 _11578_ (.A(_04050_),
    .B(_04246_),
    .Y(_04365_));
 sky130_fd_sc_hd__nor3b_1 _11579_ (.A(_04230_),
    .B(_04231_),
    .C_N(_04236_),
    .Y(_04366_));
 sky130_fd_sc_hd__a22oi_1 _11580_ (.A1(_02712_),
    .A2(_03444_),
    .B1(_05948_),
    .B2(_06682_),
    .Y(_04367_));
 sky130_fd_sc_hd__and4_1 _11581_ (.A(_02658_),
    .B(net39),
    .C(_03082_),
    .D(_00789_),
    .X(_04368_));
 sky130_fd_sc_hd__or2_1 _11582_ (.A(_04367_),
    .B(_04368_),
    .X(_04370_));
 sky130_fd_sc_hd__a21o_1 _11583_ (.A1(_04225_),
    .A2(_04226_),
    .B1(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__nand3_1 _11584_ (.A(_04225_),
    .B(_04226_),
    .C(_04370_),
    .Y(_04372_));
 sky130_fd_sc_hd__and2_1 _11585_ (.A(_04371_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__a22oi_1 _11586_ (.A1(_00878_),
    .A2(_05767_),
    .B1(_03257_),
    .B2(_00877_),
    .Y(_04374_));
 sky130_fd_sc_hd__and4_1 _11587_ (.A(_02754_),
    .B(_02797_),
    .C(_00385_),
    .D(_00783_),
    .X(_04375_));
 sky130_fd_sc_hd__nor2_1 _11588_ (.A(_04374_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand2_1 _11589_ (.A(_06608_),
    .B(_03449_),
    .Y(_04377_));
 sky130_fd_sc_hd__xnor2_1 _11590_ (.A(_04376_),
    .B(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__xor2_1 _11591_ (.A(_04373_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__o21a_1 _11592_ (.A1(_04230_),
    .A2(_04366_),
    .B1(_04379_),
    .X(_04381_));
 sky130_fd_sc_hd__nor3_1 _11593_ (.A(_04230_),
    .B(_04366_),
    .C(_04379_),
    .Y(_04382_));
 sky130_fd_sc_hd__or2_1 _11594_ (.A(_04381_),
    .B(_04382_),
    .X(_04383_));
 sky130_fd_sc_hd__inv_2 _11595_ (.A(_04219_),
    .Y(_04384_));
 sky130_fd_sc_hd__and3_1 _11596_ (.A(_04239_),
    .B(_04237_),
    .C(_04238_),
    .X(_04385_));
 sky130_fd_sc_hd__o21bai_1 _11597_ (.A1(_04232_),
    .A2(_04235_),
    .B1_N(_04233_),
    .Y(_04386_));
 sky130_fd_sc_hd__a22o_1 _11598_ (.A1(_00046_),
    .A2(_03424_),
    .B1(_03425_),
    .B2(_00049_),
    .X(_04387_));
 sky130_fd_sc_hd__nand4_1 _11599_ (.A(_00063_),
    .B(_00216_),
    .C(_05574_),
    .D(_03425_),
    .Y(_04388_));
 sky130_fd_sc_hd__a22o_1 _11600_ (.A1(_00444_),
    .A2(_05520_),
    .B1(_04387_),
    .B2(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__nand4_1 _11601_ (.A(_00221_),
    .B(_05520_),
    .C(_04387_),
    .D(_04388_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand3_1 _11602_ (.A(_04386_),
    .B(_04389_),
    .C(_04390_),
    .Y(_04392_));
 sky130_fd_sc_hd__a21o_1 _11603_ (.A1(_04389_),
    .A2(_04390_),
    .B1(_04386_),
    .X(_04393_));
 sky130_fd_sc_hd__nand2_1 _11604_ (.A(_04190_),
    .B(_04192_),
    .Y(_04394_));
 sky130_fd_sc_hd__a21o_1 _11605_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04394_),
    .X(_04395_));
 sky130_fd_sc_hd__nand3_1 _11606_ (.A(_04394_),
    .B(_04392_),
    .C(_04393_),
    .Y(_04396_));
 sky130_fd_sc_hd__a21bo_1 _11607_ (.A1(_04195_),
    .A2(_04194_),
    .B1_N(_04193_),
    .X(_04397_));
 sky130_fd_sc_hd__nand3_2 _11608_ (.A(_04395_),
    .B(_04396_),
    .C(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a21o_1 _11609_ (.A1(_04395_),
    .A2(_04396_),
    .B1(_04397_),
    .X(_04399_));
 sky130_fd_sc_hd__a22oi_1 _11610_ (.A1(_01146_),
    .A2(_00002_),
    .B1(_06561_),
    .B2(_01147_),
    .Y(_04400_));
 sky130_fd_sc_hd__and4_1 _11611_ (.A(_00124_),
    .B(_00125_),
    .C(_06525_),
    .D(_05252_),
    .X(_04401_));
 sky130_fd_sc_hd__nor2_1 _11612_ (.A(_04400_),
    .B(_04401_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _11613_ (.A(_00270_),
    .B(_00423_),
    .Y(_04404_));
 sky130_fd_sc_hd__xnor2_1 _11614_ (.A(_04403_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__a22oi_2 _11615_ (.A1(_00132_),
    .A2(_00530_),
    .B1(_05445_),
    .B2(_00133_),
    .Y(_04406_));
 sky130_fd_sc_hd__and4_1 _11616_ (.A(_00086_),
    .B(_00081_),
    .C(_06476_),
    .D(_06489_),
    .X(_04407_));
 sky130_fd_sc_hd__nand2_1 _11617_ (.A(_00088_),
    .B(_03047_),
    .Y(_04408_));
 sky130_fd_sc_hd__or3_1 _11618_ (.A(_04406_),
    .B(_04407_),
    .C(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__o21ai_1 _11619_ (.A1(_04406_),
    .A2(_04407_),
    .B1(_04408_),
    .Y(_04410_));
 sky130_fd_sc_hd__a22o_1 _11620_ (.A1(_00132_),
    .A2(_05316_),
    .B1(_05380_),
    .B2(_00133_),
    .X(_04411_));
 sky130_fd_sc_hd__a31o_1 _11621_ (.A1(_00262_),
    .A2(_05262_),
    .A3(_04411_),
    .B1(_04210_),
    .X(_04412_));
 sky130_fd_sc_hd__and3_1 _11622_ (.A(_04409_),
    .B(_04410_),
    .C(_04412_),
    .X(_04414_));
 sky130_fd_sc_hd__a21o_1 _11623_ (.A1(_04409_),
    .A2(_04410_),
    .B1(_04412_),
    .X(_04415_));
 sky130_fd_sc_hd__and2b_1 _11624_ (.A_N(_04414_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__xor2_1 _11625_ (.A(_04405_),
    .B(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__a21o_1 _11626_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__nand3_2 _11627_ (.A(_04417_),
    .B(_04398_),
    .C(_04399_),
    .Y(_04419_));
 sky130_fd_sc_hd__o211a_2 _11628_ (.A1(_04385_),
    .A2(_04244_),
    .B1(_04418_),
    .C1(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__a211oi_2 _11629_ (.A1(_04418_),
    .A2(_04419_),
    .B1(_04385_),
    .C1(_04244_),
    .Y(_04421_));
 sky130_fd_sc_hd__a211oi_4 _11630_ (.A1(_04200_),
    .A2(_04384_),
    .B1(_04420_),
    .C1(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__o211a_1 _11631_ (.A1(_04420_),
    .A2(_04421_),
    .B1(_04200_),
    .C1(_04384_),
    .X(_04423_));
 sky130_fd_sc_hd__or3_1 _11632_ (.A(_04383_),
    .B(_04422_),
    .C(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__o21ai_2 _11633_ (.A1(_04422_),
    .A2(_04423_),
    .B1(_04383_),
    .Y(_04425_));
 sky130_fd_sc_hd__o211ai_4 _11634_ (.A1(_04365_),
    .A2(_04249_),
    .B1(_04424_),
    .C1(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a211o_1 _11635_ (.A1(_04424_),
    .A2(_04425_),
    .B1(_04365_),
    .C1(_04249_),
    .X(_04427_));
 sky130_fd_sc_hd__inv_2 _11636_ (.A(_04287_),
    .Y(_04428_));
 sky130_fd_sc_hd__and3_1 _11637_ (.A(_04269_),
    .B(_04287_),
    .C(_04288_),
    .X(_04429_));
 sky130_fd_sc_hd__a211o_1 _11638_ (.A1(_04045_),
    .A2(_04048_),
    .B1(_04218_),
    .C1(_04219_),
    .X(_04430_));
 sky130_fd_sc_hd__and3_1 _11639_ (.A(_06434_),
    .B(_03604_),
    .C(_06612_),
    .X(_04431_));
 sky130_fd_sc_hd__a22o_1 _11640_ (.A1(_03604_),
    .A2(_06612_),
    .B1(_06603_),
    .B2(_06434_),
    .X(_04432_));
 sky130_fd_sc_hd__a21bo_1 _11641_ (.A1(_00445_),
    .A2(_04431_),
    .B1_N(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__nand2_1 _11642_ (.A(_02965_),
    .B(_04725_),
    .Y(_04435_));
 sky130_fd_sc_hd__xor2_4 _11643_ (.A(_04433_),
    .B(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__a32o_2 _11644_ (.A1(_03525_),
    .A2(_04660_),
    .A3(_04256_),
    .B1(_04255_),
    .B2(_04800_),
    .X(_04437_));
 sky130_fd_sc_hd__xor2_4 _11645_ (.A(_04436_),
    .B(_04437_),
    .X(_04438_));
 sky130_fd_sc_hd__and2_2 _11646_ (.A(_03722_),
    .B(_04660_),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_4 _11647_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__and2_1 _11648_ (.A(_04259_),
    .B(_04260_),
    .X(_04441_));
 sky130_fd_sc_hd__a21oi_2 _11649_ (.A1(_04261_),
    .A2(_04263_),
    .B1(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__xor2_4 _11650_ (.A(_04440_),
    .B(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__nand2_1 _11651_ (.A(_00502_),
    .B(_04607_),
    .Y(_04444_));
 sky130_fd_sc_hd__xnor2_4 _11652_ (.A(_04443_),
    .B(_04444_),
    .Y(_04446_));
 sky130_fd_sc_hd__a211oi_2 _11653_ (.A1(_04121_),
    .A2(_04126_),
    .B1(_04283_),
    .C1(_04284_),
    .Y(_04447_));
 sky130_fd_sc_hd__a21o_1 _11654_ (.A1(_04206_),
    .A2(_04215_),
    .B1(_04214_),
    .X(_04448_));
 sky130_fd_sc_hd__o21bai_1 _11655_ (.A1(_04202_),
    .A2(_04205_),
    .B1_N(_04203_),
    .Y(_04449_));
 sky130_fd_sc_hd__a22o_1 _11656_ (.A1(_02980_),
    .A2(_04972_),
    .B1(_05036_),
    .B2(_00281_),
    .X(_04450_));
 sky130_fd_sc_hd__nand4_1 _11657_ (.A(_02983_),
    .B(_02984_),
    .C(_04972_),
    .D(_00421_),
    .Y(_04451_));
 sky130_fd_sc_hd__a22o_1 _11658_ (.A1(_00345_),
    .A2(_04918_),
    .B1(_04450_),
    .B2(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__nand4_1 _11659_ (.A(_02987_),
    .B(_04918_),
    .C(_04450_),
    .D(_04451_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_1 _11660_ (.A(_04449_),
    .B(_04452_),
    .C(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21o_1 _11661_ (.A1(_04452_),
    .A2(_04453_),
    .B1(_04449_),
    .X(_04455_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_04275_),
    .B(_04277_),
    .Y(_04457_));
 sky130_fd_sc_hd__a21o_1 _11663_ (.A1(_04454_),
    .A2(_04455_),
    .B1(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__nand3_1 _11664_ (.A(_04457_),
    .B(_04454_),
    .C(_04455_),
    .Y(_04459_));
 sky130_fd_sc_hd__and3_2 _11665_ (.A(_04448_),
    .B(_04458_),
    .C(_04459_),
    .X(_04460_));
 sky130_fd_sc_hd__a21oi_1 _11666_ (.A1(_04458_),
    .A2(_04459_),
    .B1(_04448_),
    .Y(_04461_));
 sky130_fd_sc_hd__a211o_1 _11667_ (.A1(_04278_),
    .A2(_04282_),
    .B1(_04460_),
    .C1(_04461_),
    .X(_04462_));
 sky130_fd_sc_hd__o211ai_1 _11668_ (.A1(_04460_),
    .A2(_04461_),
    .B1(_04278_),
    .C1(_04282_),
    .Y(_04463_));
 sky130_fd_sc_hd__o211ai_2 _11669_ (.A1(_04283_),
    .A2(_04447_),
    .B1(_04462_),
    .C1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__a211o_1 _11670_ (.A1(_04462_),
    .A2(_04463_),
    .B1(_04283_),
    .C1(_04447_),
    .X(_04465_));
 sky130_fd_sc_hd__and3_2 _11671_ (.A(_04446_),
    .B(_04464_),
    .C(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__a21oi_1 _11672_ (.A1(_04464_),
    .A2(_04465_),
    .B1(_04446_),
    .Y(_04468_));
 sky130_fd_sc_hd__a211o_2 _11673_ (.A1(_04430_),
    .A2(_04222_),
    .B1(_04466_),
    .C1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o211ai_2 _11674_ (.A1(_04466_),
    .A2(_04468_),
    .B1(_04430_),
    .C1(_04222_),
    .Y(_04470_));
 sky130_fd_sc_hd__o211ai_4 _11675_ (.A1(_04428_),
    .A2(_04429_),
    .B1(_04469_),
    .C1(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__a211o_1 _11676_ (.A1(_04469_),
    .A2(_04470_),
    .B1(_04428_),
    .C1(_04429_),
    .X(_04472_));
 sky130_fd_sc_hd__and4_1 _11677_ (.A(_04426_),
    .B(_04427_),
    .C(_04471_),
    .D(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__a22oi_2 _11678_ (.A1(_04426_),
    .A2(_04427_),
    .B1(_04471_),
    .B2(_04472_),
    .Y(_04474_));
 sky130_fd_sc_hd__a211oi_4 _11679_ (.A1(_04250_),
    .A2(_04364_),
    .B1(_04473_),
    .C1(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__o211a_1 _11680_ (.A1(_04473_),
    .A2(_04474_),
    .B1(_04250_),
    .C1(_04364_),
    .X(_04476_));
 sky130_fd_sc_hd__a211o_1 _11681_ (.A1(_04291_),
    .A2(_04293_),
    .B1(_04475_),
    .C1(_04476_),
    .X(_04477_));
 sky130_fd_sc_hd__o211ai_2 _11682_ (.A1(_04475_),
    .A2(_04476_),
    .B1(_04291_),
    .C1(_04293_),
    .Y(_04479_));
 sky130_fd_sc_hd__o211a_2 _11683_ (.A1(_04298_),
    .A2(_04363_),
    .B1(_04477_),
    .C1(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__a211oi_4 _11684_ (.A1(_04477_),
    .A2(_04479_),
    .B1(_04298_),
    .C1(_04363_),
    .Y(_04481_));
 sky130_fd_sc_hd__a211oi_1 _11685_ (.A1(_04361_),
    .A2(_04362_),
    .B1(_04480_),
    .C1(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__o211a_1 _11686_ (.A1(_04480_),
    .A2(_04481_),
    .B1(_04361_),
    .C1(_04362_),
    .X(_04483_));
 sky130_fd_sc_hd__a211o_1 _11687_ (.A1(_04360_),
    .A2(_04304_),
    .B1(_04482_),
    .C1(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__inv_2 _11688_ (.A(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__o211a_1 _11689_ (.A1(_04482_),
    .A2(_04483_),
    .B1(_04360_),
    .C1(_04304_),
    .X(_04486_));
 sky130_fd_sc_hd__nor2_1 _11690_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__a21oi_1 _11691_ (.A1(_04359_),
    .A2(_04487_),
    .B1(_06428_),
    .Y(_04488_));
 sky130_fd_sc_hd__o21ai_1 _11692_ (.A1(_04359_),
    .A2(_04487_),
    .B1(_04488_),
    .Y(_04490_));
 sky130_fd_sc_hd__o311a_1 _11693_ (.A1(_02571_),
    .A2(_04159_),
    .A3(_04348_),
    .B1(_04357_),
    .C1(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__o21ai_4 _11694_ (.A1(_02713_),
    .A2(_04346_),
    .B1(_04491_),
    .Y(net100));
 sky130_fd_sc_hd__or2b_1 _11695_ (.A(_02789_),
    .B_N(_02785_),
    .X(_04492_));
 sky130_fd_sc_hd__o211a_1 _11696_ (.A1(_02791_),
    .A2(_04343_),
    .B1(_04492_),
    .C1(_02787_),
    .X(_04493_));
 sky130_fd_sc_hd__mux2_1 _11697_ (.A0(_04493_),
    .A1(_02891_),
    .S(_02928_),
    .X(_04494_));
 sky130_fd_sc_hd__or2_1 _11698_ (.A(_02860_),
    .B(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__nand2_1 _11699_ (.A(_02860_),
    .B(_04494_),
    .Y(_04496_));
 sky130_fd_sc_hd__a211oi_2 _11700_ (.A1(_04291_),
    .A2(_04293_),
    .B1(_04475_),
    .C1(_04476_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand4_1 _11701_ (.A(_04426_),
    .B(_04427_),
    .C(_04471_),
    .D(_04472_),
    .Y(_04498_));
 sky130_fd_sc_hd__nor3_1 _11702_ (.A(_04383_),
    .B(_04422_),
    .C(_04423_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _11703_ (.A(_04373_),
    .B(_04378_),
    .Y(_04500_));
 sky130_fd_sc_hd__and3_1 _11704_ (.A(_00877_),
    .B(_00878_),
    .C(_05820_),
    .X(_04501_));
 sky130_fd_sc_hd__a22o_1 _11705_ (.A1(_00878_),
    .A2(_05820_),
    .B1(_03444_),
    .B2(_00012_),
    .X(_04502_));
 sky130_fd_sc_hd__a21bo_1 _11706_ (.A1(_05895_),
    .A2(_04501_),
    .B1_N(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__nand2_1 _11707_ (.A(_02851_),
    .B(_05777_),
    .Y(_04504_));
 sky130_fd_sc_hd__xor2_1 _11708_ (.A(_04503_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__nand2_1 _11709_ (.A(_02669_),
    .B(_05906_),
    .Y(_04506_));
 sky130_fd_sc_hd__and3_1 _11710_ (.A(_02723_),
    .B(_05970_),
    .C(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__xnor2_1 _11711_ (.A(_04505_),
    .B(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21oi_1 _11712_ (.A1(_04371_),
    .A2(_04500_),
    .B1(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__and3_1 _11713_ (.A(_04371_),
    .B(_04500_),
    .C(_04508_),
    .X(_04511_));
 sky130_fd_sc_hd__or2_1 _11714_ (.A(_04510_),
    .B(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__o21bai_1 _11715_ (.A1(_04374_),
    .A2(_04377_),
    .B1_N(_04375_),
    .Y(_04513_));
 sky130_fd_sc_hd__a22o_1 _11716_ (.A1(_00046_),
    .A2(_00382_),
    .B1(_00163_),
    .B2(_00049_),
    .X(_04514_));
 sky130_fd_sc_hd__nand4_1 _11717_ (.A(_00063_),
    .B(_00062_),
    .C(_03425_),
    .D(_05702_),
    .Y(_04515_));
 sky130_fd_sc_hd__a22o_1 _11718_ (.A1(_00058_),
    .A2(_03071_),
    .B1(_04514_),
    .B2(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__nand4_1 _11719_ (.A(_00221_),
    .B(_05585_),
    .C(_04514_),
    .D(_04515_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand3_1 _11720_ (.A(_04513_),
    .B(_04516_),
    .C(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21o_1 _11721_ (.A1(_04516_),
    .A2(_04517_),
    .B1(_04513_),
    .X(_04519_));
 sky130_fd_sc_hd__nand2_1 _11722_ (.A(_04388_),
    .B(_04390_),
    .Y(_04521_));
 sky130_fd_sc_hd__a21o_1 _11723_ (.A1(_04518_),
    .A2(_04519_),
    .B1(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__nand3_1 _11724_ (.A(_04521_),
    .B(_04518_),
    .C(_04519_),
    .Y(_04523_));
 sky130_fd_sc_hd__a21bo_1 _11725_ (.A1(_04394_),
    .A2(_04393_),
    .B1_N(_04392_),
    .X(_04524_));
 sky130_fd_sc_hd__nand3_1 _11726_ (.A(_04522_),
    .B(_04523_),
    .C(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__a21o_1 _11727_ (.A1(_04522_),
    .A2(_04523_),
    .B1(_04524_),
    .X(_04526_));
 sky130_fd_sc_hd__a22oi_2 _11728_ (.A1(_01146_),
    .A2(_06561_),
    .B1(_03047_),
    .B2(_01147_),
    .Y(_04527_));
 sky130_fd_sc_hd__and4_1 _11729_ (.A(_00124_),
    .B(_00125_),
    .C(_05252_),
    .D(_05316_),
    .X(_04528_));
 sky130_fd_sc_hd__nand2_1 _11730_ (.A(_03324_),
    .B(_05198_),
    .Y(_04529_));
 sky130_fd_sc_hd__or3_1 _11731_ (.A(_04527_),
    .B(_04528_),
    .C(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__o21ai_1 _11732_ (.A1(_04527_),
    .A2(_04528_),
    .B1(_04529_),
    .Y(_04532_));
 sky130_fd_sc_hd__nand2_1 _11733_ (.A(_04530_),
    .B(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__a22oi_2 _11734_ (.A1(_03099_),
    .A2(_06666_),
    .B1(_00398_),
    .B2(_03056_),
    .Y(_04534_));
 sky130_fd_sc_hd__and4_1 _11735_ (.A(_00237_),
    .B(_00462_),
    .C(_06489_),
    .D(_05498_),
    .X(_04535_));
 sky130_fd_sc_hd__nand2_1 _11736_ (.A(_00088_),
    .B(_05380_),
    .Y(_04536_));
 sky130_fd_sc_hd__or3_1 _11737_ (.A(_04534_),
    .B(_04535_),
    .C(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__o21ai_1 _11738_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04536_),
    .Y(_04538_));
 sky130_fd_sc_hd__o21bai_1 _11739_ (.A1(_04406_),
    .A2(_04408_),
    .B1_N(_04407_),
    .Y(_04539_));
 sky130_fd_sc_hd__and3_1 _11740_ (.A(_04537_),
    .B(_04538_),
    .C(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__a21oi_1 _11741_ (.A1(_04537_),
    .A2(_04538_),
    .B1(_04539_),
    .Y(_04541_));
 sky130_fd_sc_hd__nor2_1 _11742_ (.A(_04540_),
    .B(_04541_),
    .Y(_04543_));
 sky130_fd_sc_hd__xnor2_1 _11743_ (.A(_04533_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__a21o_1 _11744_ (.A1(_04525_),
    .A2(_04526_),
    .B1(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__nand3_1 _11745_ (.A(_04544_),
    .B(_04525_),
    .C(_04526_),
    .Y(_04546_));
 sky130_fd_sc_hd__and3_1 _11746_ (.A(_04381_),
    .B(_04545_),
    .C(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__a21oi_1 _11747_ (.A1(_04545_),
    .A2(_04546_),
    .B1(_04381_),
    .Y(_04548_));
 sky130_fd_sc_hd__a211oi_2 _11748_ (.A1(_04398_),
    .A2(_04419_),
    .B1(_04547_),
    .C1(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__o211a_1 _11749_ (.A1(_04547_),
    .A2(_04548_),
    .B1(_04398_),
    .C1(_04419_),
    .X(_04550_));
 sky130_fd_sc_hd__or3_1 _11750_ (.A(_04512_),
    .B(_04549_),
    .C(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__o21ai_1 _11751_ (.A1(_04549_),
    .A2(_04550_),
    .B1(_04512_),
    .Y(_04552_));
 sky130_fd_sc_hd__and3_1 _11752_ (.A(_04499_),
    .B(_04551_),
    .C(_04552_),
    .X(_04554_));
 sky130_fd_sc_hd__a21oi_1 _11753_ (.A1(_04551_),
    .A2(_04552_),
    .B1(_04499_),
    .Y(_04555_));
 sky130_fd_sc_hd__inv_2 _11754_ (.A(_04464_),
    .Y(_04556_));
 sky130_fd_sc_hd__and3_1 _11755_ (.A(_03539_),
    .B(_00678_),
    .C(_06603_),
    .X(_04557_));
 sky130_fd_sc_hd__a22o_1 _11756_ (.A1(_00678_),
    .A2(_06603_),
    .B1(_06605_),
    .B2(_03539_),
    .X(_04558_));
 sky130_fd_sc_hd__a21bo_2 _11757_ (.A1(_00550_),
    .A2(_04557_),
    .B1_N(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_03658_),
    .B(_06613_),
    .Y(_04560_));
 sky130_fd_sc_hd__xor2_4 _11759_ (.A(_04559_),
    .B(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__a32o_2 _11760_ (.A1(_03525_),
    .A2(_04725_),
    .A3(_04432_),
    .B1(_04431_),
    .B2(_04854_),
    .X(_04562_));
 sky130_fd_sc_hd__xor2_4 _11761_ (.A(_04561_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_06429_),
    .B(_04725_),
    .Y(_04564_));
 sky130_fd_sc_hd__xor2_4 _11763_ (.A(_04563_),
    .B(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__and2_1 _11764_ (.A(_04436_),
    .B(_04437_),
    .X(_04566_));
 sky130_fd_sc_hd__a21oi_2 _11765_ (.A1(_04438_),
    .A2(_04439_),
    .B1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__xor2_4 _11766_ (.A(_04565_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_00502_),
    .B(_04660_),
    .Y(_04569_));
 sky130_fd_sc_hd__xnor2_4 _11768_ (.A(_04568_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__a211oi_2 _11769_ (.A1(_04278_),
    .A2(_04282_),
    .B1(_04460_),
    .C1(_04461_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21o_1 _11770_ (.A1(_04405_),
    .A2(_04415_),
    .B1(_04414_),
    .X(_04572_));
 sky130_fd_sc_hd__o21bai_1 _11771_ (.A1(_04400_),
    .A2(_04404_),
    .B1_N(_04401_),
    .Y(_04573_));
 sky130_fd_sc_hd__a22o_1 _11772_ (.A1(_00289_),
    .A2(_05036_),
    .B1(_05112_),
    .B2(_00290_),
    .X(_04575_));
 sky130_fd_sc_hd__nand4_2 _11773_ (.A(_00281_),
    .B(_03443_),
    .C(_05036_),
    .D(_00534_),
    .Y(_04576_));
 sky130_fd_sc_hd__a22o_1 _11774_ (.A1(_00283_),
    .A2(_00197_),
    .B1(_04575_),
    .B2(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__nand4_2 _11775_ (.A(_00345_),
    .B(_00197_),
    .C(_04575_),
    .D(_04576_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand3_2 _11776_ (.A(_04573_),
    .B(_04577_),
    .C(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__a21o_1 _11777_ (.A1(_04577_),
    .A2(_04578_),
    .B1(_04573_),
    .X(_04580_));
 sky130_fd_sc_hd__nand2_1 _11778_ (.A(_04451_),
    .B(_04453_),
    .Y(_04581_));
 sky130_fd_sc_hd__a21o_1 _11779_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_04581_),
    .X(_04582_));
 sky130_fd_sc_hd__nand3_2 _11780_ (.A(_04581_),
    .B(_04579_),
    .C(_04580_),
    .Y(_04583_));
 sky130_fd_sc_hd__and3_1 _11781_ (.A(_04572_),
    .B(_04582_),
    .C(_04583_),
    .X(_04584_));
 sky130_fd_sc_hd__a21oi_1 _11782_ (.A1(_04582_),
    .A2(_04583_),
    .B1(_04572_),
    .Y(_04586_));
 sky130_fd_sc_hd__a211o_1 _11783_ (.A1(_04454_),
    .A2(_04459_),
    .B1(_04584_),
    .C1(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__o211ai_1 _11784_ (.A1(_04584_),
    .A2(_04586_),
    .B1(_04454_),
    .C1(_04459_),
    .Y(_04588_));
 sky130_fd_sc_hd__o211ai_2 _11785_ (.A1(_04460_),
    .A2(_04571_),
    .B1(_04587_),
    .C1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__a211o_1 _11786_ (.A1(_04587_),
    .A2(_04588_),
    .B1(_04460_),
    .C1(_04571_),
    .X(_04590_));
 sky130_fd_sc_hd__nand3_2 _11787_ (.A(_04570_),
    .B(_04589_),
    .C(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a21o_1 _11788_ (.A1(_04589_),
    .A2(_04590_),
    .B1(_04570_),
    .X(_04592_));
 sky130_fd_sc_hd__o211ai_4 _11789_ (.A1(_04420_),
    .A2(_04422_),
    .B1(_04591_),
    .C1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__a211o_1 _11790_ (.A1(_04591_),
    .A2(_04592_),
    .B1(_04420_),
    .C1(_04422_),
    .X(_04594_));
 sky130_fd_sc_hd__o211ai_4 _11791_ (.A1(_04556_),
    .A2(_04466_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__a211o_1 _11792_ (.A1(_04593_),
    .A2(_04594_),
    .B1(_04556_),
    .C1(_04466_),
    .X(_04597_));
 sky130_fd_sc_hd__and4bb_1 _11793_ (.A_N(_04554_),
    .B_N(_04555_),
    .C(_04595_),
    .D(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__a2bb2oi_1 _11794_ (.A1_N(_04554_),
    .A2_N(_04555_),
    .B1(_04595_),
    .B2(_04597_),
    .Y(_04599_));
 sky130_fd_sc_hd__a211oi_1 _11795_ (.A1(_04426_),
    .A2(_04498_),
    .B1(_04598_),
    .C1(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__o211a_1 _11796_ (.A1(_04598_),
    .A2(_04599_),
    .B1(_04426_),
    .C1(_04498_),
    .X(_04601_));
 sky130_fd_sc_hd__a211o_2 _11797_ (.A1(_04469_),
    .A2(_04471_),
    .B1(_04600_),
    .C1(_04601_),
    .X(_04602_));
 sky130_fd_sc_hd__o211ai_2 _11798_ (.A1(_04600_),
    .A2(_04601_),
    .B1(_04469_),
    .C1(_04471_),
    .Y(_04603_));
 sky130_fd_sc_hd__o211ai_4 _11799_ (.A1(_04475_),
    .A2(_04497_),
    .B1(_04602_),
    .C1(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__a211o_1 _11800_ (.A1(_04602_),
    .A2(_04603_),
    .B1(_04475_),
    .C1(_04497_),
    .X(_04605_));
 sky130_fd_sc_hd__and2_2 _11801_ (.A(_04604_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__nor2_1 _11802_ (.A(_04440_),
    .B(_04442_),
    .Y(_04608_));
 sky130_fd_sc_hd__a31o_1 _11803_ (.A1(_03820_),
    .A2(_04607_),
    .A3(_04443_),
    .B1(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__nand2_1 _11804_ (.A(_04606_),
    .B(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__or2_1 _11805_ (.A(_04606_),
    .B(_04609_),
    .X(_04611_));
 sky130_fd_sc_hd__nand2_1 _11806_ (.A(_04610_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _11807_ (.A(_04480_),
    .B(_04482_),
    .Y(_04613_));
 sky130_fd_sc_hd__xnor2_1 _11808_ (.A(_04612_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _11809_ (.A(_04312_),
    .B(_04487_),
    .Y(_04615_));
 sky130_fd_sc_hd__a21o_1 _11810_ (.A1(_04310_),
    .A2(_04484_),
    .B1(_04486_),
    .X(_04616_));
 sky130_fd_sc_hd__o21a_1 _11811_ (.A1(_04322_),
    .A2(_04615_),
    .B1(_04616_),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_1 _11812_ (.A(_04614_),
    .B(_04617_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor2_1 _11813_ (.A(_04614_),
    .B(_04617_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _11814_ (.A(_06428_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__or2b_1 _11815_ (.A(_02572_),
    .B_N(_02551_),
    .X(_04622_));
 sky130_fd_sc_hd__xnor2_1 _11816_ (.A(_04622_),
    .B(_02571_),
    .Y(_04623_));
 sky130_fd_sc_hd__o21a_1 _11817_ (.A1(_02790_),
    .A2(_04349_),
    .B1(_01350_),
    .X(_04624_));
 sky130_fd_sc_hd__xnor2_1 _11818_ (.A(_02860_),
    .B(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__a2bb2o_1 _11819_ (.A1_N(_04607_),
    .A2_N(_02941_),
    .B1(_02731_),
    .B2(\AuI.result[10] ),
    .X(_04626_));
 sky130_fd_sc_hd__buf_2 _11820_ (.A(_06045_),
    .X(_04627_));
 sky130_fd_sc_hd__a32o_1 _11821_ (.A1(_02669_),
    .A2(_04607_),
    .A3(_02743_),
    .B1(_02944_),
    .B2(_04542_),
    .X(_04628_));
 sky130_fd_sc_hd__a221o_1 _11822_ (.A1(\MuI.result[10] ),
    .A2(_02737_),
    .B1(_04011_),
    .B2(_02860_),
    .C1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__a221o_1 _11823_ (.A1(\FuI.Integer[10] ),
    .A2(_04627_),
    .B1(_03675_),
    .B2(_04671_),
    .C1(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__a211o_1 _11824_ (.A1(_02669_),
    .A2(_02724_),
    .B1(_04626_),
    .C1(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__a21o_1 _11825_ (.A1(_03489_),
    .A2(_04625_),
    .B1(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__a221o_1 _11826_ (.A1(_04619_),
    .A2(_04621_),
    .B1(_04623_),
    .B2(_03315_),
    .C1(_04632_),
    .X(_04633_));
 sky130_fd_sc_hd__a31o_2 _11827_ (.A1(_02752_),
    .A2(_04495_),
    .A3(_04496_),
    .B1(_04633_),
    .X(net70));
 sky130_fd_sc_hd__o21ai_1 _11828_ (.A1(_02860_),
    .A2(_04493_),
    .B1(_02858_),
    .Y(_04634_));
 sky130_fd_sc_hd__buf_4 _11829_ (.A(_02926_),
    .X(_04635_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(_04634_),
    .A1(_02892_),
    .S(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(_02871_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__or2_1 _11832_ (.A(_02871_),
    .B(_04636_),
    .X(_04639_));
 sky130_fd_sc_hd__or2b_1 _11833_ (.A(_02574_),
    .B_N(_02521_),
    .X(_04640_));
 sky130_fd_sc_hd__xnor2_1 _11834_ (.A(_04640_),
    .B(_02573_),
    .Y(_04641_));
 sky130_fd_sc_hd__clkbuf_4 _11835_ (.A(_02944_),
    .X(_04642_));
 sky130_fd_sc_hd__o22ai_1 _11836_ (.A1(_04671_),
    .A2(_02941_),
    .B1(_02871_),
    .B2(_03306_),
    .Y(_04643_));
 sky130_fd_sc_hd__a221o_1 _11837_ (.A1(\MuI.result[11] ),
    .A2(_02738_),
    .B1(_04642_),
    .B2(_04607_),
    .C1(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__a32o_1 _11838_ (.A1(_02723_),
    .A2(_04671_),
    .A3(_02744_),
    .B1(_04627_),
    .B2(\FuI.Integer[11] ),
    .X(_04645_));
 sky130_fd_sc_hd__a221o_1 _11839_ (.A1(_04736_),
    .A2(_02719_),
    .B1(_02722_),
    .B2(_02723_),
    .C1(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__o21a_1 _11840_ (.A1(_02861_),
    .A2(_04624_),
    .B1(_01349_),
    .X(_04647_));
 sky130_fd_sc_hd__xor2_1 _11841_ (.A(_02871_),
    .B(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__a22o_1 _11842_ (.A1(\AuI.result[11] ),
    .A2(_02732_),
    .B1(_04648_),
    .B2(_02935_),
    .X(_04650_));
 sky130_fd_sc_hd__or3_1 _11843_ (.A(_04644_),
    .B(_04646_),
    .C(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__or2_1 _11844_ (.A(_04565_),
    .B(_04567_),
    .X(_04652_));
 sky130_fd_sc_hd__nand3_1 _11845_ (.A(_03831_),
    .B(_04671_),
    .C(_04568_),
    .Y(_04653_));
 sky130_fd_sc_hd__a211o_1 _11846_ (.A1(_04426_),
    .A2(_04498_),
    .B1(_04598_),
    .C1(_04599_),
    .X(_04654_));
 sky130_fd_sc_hd__and3_1 _11847_ (.A(_00877_),
    .B(_00011_),
    .C(_03444_),
    .X(_04655_));
 sky130_fd_sc_hd__a22o_1 _11848_ (.A1(_00878_),
    .A2(_03444_),
    .B1(_05948_),
    .B2(_00012_),
    .X(_04656_));
 sky130_fd_sc_hd__a21bo_1 _11849_ (.A1(_05970_),
    .A2(_04655_),
    .B1_N(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _11850_ (.A(_02862_),
    .B(_05831_),
    .Y(_04658_));
 sky130_fd_sc_hd__xor2_1 _11851_ (.A(_04657_),
    .B(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__a21oi_1 _11852_ (.A1(_04505_),
    .A2(_04507_),
    .B1(_04368_),
    .Y(_04661_));
 sky130_fd_sc_hd__xnor2_1 _11853_ (.A(_04659_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__a32o_1 _11854_ (.A1(_06610_),
    .A2(_05777_),
    .A3(_04502_),
    .B1(_04501_),
    .B2(_05895_),
    .X(_04663_));
 sky130_fd_sc_hd__a22o_1 _11855_ (.A1(_00216_),
    .A2(_05702_),
    .B1(_05767_),
    .B2(_00217_),
    .X(_04664_));
 sky130_fd_sc_hd__nand4_1 _11856_ (.A(_02905_),
    .B(_02959_),
    .C(_03449_),
    .D(_05767_),
    .Y(_04665_));
 sky130_fd_sc_hd__a22o_1 _11857_ (.A1(_00221_),
    .A2(_05660_),
    .B1(_04664_),
    .B2(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__nand4_1 _11858_ (.A(_03013_),
    .B(_05660_),
    .C(_04664_),
    .D(_04665_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand3_1 _11859_ (.A(_04663_),
    .B(_04666_),
    .C(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__a21o_1 _11860_ (.A1(_04666_),
    .A2(_04667_),
    .B1(_04663_),
    .X(_04669_));
 sky130_fd_sc_hd__nand2_1 _11861_ (.A(_04515_),
    .B(_04517_),
    .Y(_04670_));
 sky130_fd_sc_hd__a21o_1 _11862_ (.A1(_04668_),
    .A2(_04669_),
    .B1(_04670_),
    .X(_04672_));
 sky130_fd_sc_hd__nand3_1 _11863_ (.A(_04670_),
    .B(_04668_),
    .C(_04669_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_1 _11864_ (.A(_04518_),
    .B(_04523_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand3_1 _11865_ (.A(_04672_),
    .B(_04673_),
    .C(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__a21o_1 _11866_ (.A1(_04672_),
    .A2(_04673_),
    .B1(_04674_),
    .X(_04676_));
 sky130_fd_sc_hd__nand2_2 _11867_ (.A(_00124_),
    .B(_05316_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_2 _11868_ (.A(_00125_),
    .B(_00530_),
    .Y(_04678_));
 sky130_fd_sc_hd__a22o_1 _11869_ (.A1(_03271_),
    .A2(_06562_),
    .B1(_00530_),
    .B2(_03217_),
    .X(_04679_));
 sky130_fd_sc_hd__o21a_1 _11870_ (.A1(_04677_),
    .A2(_04678_),
    .B1(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__nand2_1 _11871_ (.A(_03324_),
    .B(_05262_),
    .Y(_04681_));
 sky130_fd_sc_hd__xnor2_1 _11872_ (.A(_04680_),
    .B(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__a22oi_2 _11873_ (.A1(_00462_),
    .A2(_05498_),
    .B1(_05563_),
    .B2(_00237_),
    .Y(_04684_));
 sky130_fd_sc_hd__and4_1 _11874_ (.A(_00095_),
    .B(net117),
    .C(_06466_),
    .D(_06461_),
    .X(_04685_));
 sky130_fd_sc_hd__nand2_1 _11875_ (.A(_03152_),
    .B(_06666_),
    .Y(_04686_));
 sky130_fd_sc_hd__or3_1 _11876_ (.A(_04684_),
    .B(_04685_),
    .C(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__o21ai_1 _11877_ (.A1(_04684_),
    .A2(_04685_),
    .B1(_04686_),
    .Y(_04688_));
 sky130_fd_sc_hd__o21bai_1 _11878_ (.A1(_04534_),
    .A2(_04536_),
    .B1_N(_04535_),
    .Y(_04689_));
 sky130_fd_sc_hd__and3_1 _11879_ (.A(_04687_),
    .B(_04688_),
    .C(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__a21o_1 _11880_ (.A1(_04687_),
    .A2(_04688_),
    .B1(_04689_),
    .X(_04691_));
 sky130_fd_sc_hd__and2b_1 _11881_ (.A_N(_04690_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__xor2_1 _11882_ (.A(_04683_),
    .B(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__a21o_1 _11883_ (.A1(_04675_),
    .A2(_04676_),
    .B1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__nand3_1 _11884_ (.A(_04693_),
    .B(_04675_),
    .C(_04676_),
    .Y(_04695_));
 sky130_fd_sc_hd__and3_1 _11885_ (.A(_04510_),
    .B(_04694_),
    .C(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__a21oi_1 _11886_ (.A1(_04694_),
    .A2(_04695_),
    .B1(_04510_),
    .Y(_04697_));
 sky130_fd_sc_hd__a211o_1 _11887_ (.A1(_04525_),
    .A2(_04546_),
    .B1(_04696_),
    .C1(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__o211ai_1 _11888_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04525_),
    .C1(_04546_),
    .Y(_04699_));
 sky130_fd_sc_hd__and3_1 _11889_ (.A(_04662_),
    .B(_04698_),
    .C(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__a21oi_1 _11890_ (.A1(_04698_),
    .A2(_04699_),
    .B1(_04662_),
    .Y(_04701_));
 sky130_fd_sc_hd__or3_2 _11891_ (.A(_04551_),
    .B(_04700_),
    .C(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__o21ai_1 _11892_ (.A1(_04700_),
    .A2(_04701_),
    .B1(_04551_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _11893_ (.A(_04561_),
    .B(_04562_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand3_1 _11894_ (.A(_03744_),
    .B(_04725_),
    .C(_04563_),
    .Y(_04706_));
 sky130_fd_sc_hd__and3_1 _11895_ (.A(_06434_),
    .B(_03604_),
    .C(_06605_),
    .X(_04707_));
 sky130_fd_sc_hd__a22o_1 _11896_ (.A1(_03604_),
    .A2(_06605_),
    .B1(_06591_),
    .B2(_06434_),
    .X(_04708_));
 sky130_fd_sc_hd__a21bo_1 _11897_ (.A1(_00197_),
    .A2(_04707_),
    .B1_N(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__nand2_1 _11898_ (.A(_02965_),
    .B(_04854_),
    .Y(_04710_));
 sky130_fd_sc_hd__xor2_1 _11899_ (.A(_04709_),
    .B(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__a32o_1 _11900_ (.A1(_03525_),
    .A2(_06613_),
    .A3(_04558_),
    .B1(_04557_),
    .B2(_04918_),
    .X(_04712_));
 sky130_fd_sc_hd__xor2_1 _11901_ (.A(_04711_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__and2_1 _11902_ (.A(_03722_),
    .B(_04800_),
    .X(_04715_));
 sky130_fd_sc_hd__xnor2_1 _11903_ (.A(_04713_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hd__a21oi_1 _11904_ (.A1(_04705_),
    .A2(_04706_),
    .B1(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__and3_1 _11905_ (.A(_04705_),
    .B(_04706_),
    .C(_04716_),
    .X(_04718_));
 sky130_fd_sc_hd__nor2_1 _11906_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _11907_ (.A(_03798_),
    .B(_04736_),
    .Y(_04720_));
 sky130_fd_sc_hd__xnor2_2 _11908_ (.A(_04719_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand3_1 _11909_ (.A(_04572_),
    .B(_04582_),
    .C(_04583_),
    .Y(_04722_));
 sky130_fd_sc_hd__o21bai_1 _11910_ (.A1(_04533_),
    .A2(_04541_),
    .B1_N(_04540_),
    .Y(_04723_));
 sky130_fd_sc_hd__o21bai_1 _11911_ (.A1(_04527_),
    .A2(_04529_),
    .B1_N(_04528_),
    .Y(_04724_));
 sky130_fd_sc_hd__a22o_1 _11912_ (.A1(_03443_),
    .A2(_05112_),
    .B1(_06525_),
    .B2(_00290_),
    .X(_04726_));
 sky130_fd_sc_hd__nand4_1 _11913_ (.A(_00281_),
    .B(_02980_),
    .C(_00534_),
    .D(_00002_),
    .Y(_04727_));
 sky130_fd_sc_hd__a22o_1 _11914_ (.A1(_03486_),
    .A2(_05047_),
    .B1(_04726_),
    .B2(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__nand4_1 _11915_ (.A(_00345_),
    .B(_05047_),
    .C(_04726_),
    .D(_04727_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand3_1 _11916_ (.A(_04724_),
    .B(_04728_),
    .C(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__a21o_1 _11917_ (.A1(_04728_),
    .A2(_04729_),
    .B1(_04724_),
    .X(_04731_));
 sky130_fd_sc_hd__nand2_1 _11918_ (.A(_04576_),
    .B(_04578_),
    .Y(_04732_));
 sky130_fd_sc_hd__a21o_1 _11919_ (.A1(_04730_),
    .A2(_04731_),
    .B1(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__nand3_1 _11920_ (.A(_04732_),
    .B(_04730_),
    .C(_04731_),
    .Y(_04734_));
 sky130_fd_sc_hd__and3_1 _11921_ (.A(_04723_),
    .B(_04733_),
    .C(_04734_),
    .X(_04735_));
 sky130_fd_sc_hd__a21oi_1 _11922_ (.A1(_04733_),
    .A2(_04734_),
    .B1(_04723_),
    .Y(_04737_));
 sky130_fd_sc_hd__a211oi_2 _11923_ (.A1(_04579_),
    .A2(_04583_),
    .B1(_04735_),
    .C1(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__o211a_1 _11924_ (.A1(_04735_),
    .A2(_04737_),
    .B1(_04579_),
    .C1(_04583_),
    .X(_04739_));
 sky130_fd_sc_hd__a211o_1 _11925_ (.A1(_04722_),
    .A2(_04587_),
    .B1(_04738_),
    .C1(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__o211ai_1 _11926_ (.A1(_04738_),
    .A2(_04739_),
    .B1(_04722_),
    .C1(_04587_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand3_1 _11927_ (.A(_04721_),
    .B(_04740_),
    .C(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21o_1 _11928_ (.A1(_04740_),
    .A2(_04741_),
    .B1(_04721_),
    .X(_04743_));
 sky130_fd_sc_hd__o211a_1 _11929_ (.A1(_04547_),
    .A2(_04549_),
    .B1(_04742_),
    .C1(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__a211oi_1 _11930_ (.A1(_04742_),
    .A2(_04743_),
    .B1(_04547_),
    .C1(_04549_),
    .Y(_04745_));
 sky130_fd_sc_hd__a211o_1 _11931_ (.A1(_04589_),
    .A2(_04591_),
    .B1(_04744_),
    .C1(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__o211ai_1 _11932_ (.A1(_04744_),
    .A2(_04745_),
    .B1(_04589_),
    .C1(_04591_),
    .Y(_04748_));
 sky130_fd_sc_hd__nand4_2 _11933_ (.A(_04702_),
    .B(_04704_),
    .C(_04746_),
    .D(_04748_),
    .Y(_04749_));
 sky130_fd_sc_hd__a22o_1 _11934_ (.A1(_04702_),
    .A2(_04704_),
    .B1(_04746_),
    .B2(_04748_),
    .X(_04750_));
 sky130_fd_sc_hd__o211a_2 _11935_ (.A1(_04554_),
    .A2(_04598_),
    .B1(_04749_),
    .C1(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a211oi_2 _11936_ (.A1(_04749_),
    .A2(_04750_),
    .B1(_04554_),
    .C1(_04598_),
    .Y(_04752_));
 sky130_fd_sc_hd__a211oi_4 _11937_ (.A1(_04593_),
    .A2(_04595_),
    .B1(_04751_),
    .C1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__o211a_1 _11938_ (.A1(_04751_),
    .A2(_04752_),
    .B1(_04593_),
    .C1(_04595_),
    .X(_04754_));
 sky130_fd_sc_hd__a211oi_4 _11939_ (.A1(_04654_),
    .A2(_04602_),
    .B1(_04753_),
    .C1(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__o211a_2 _11940_ (.A1(_04753_),
    .A2(_04754_),
    .B1(_04654_),
    .C1(_04602_),
    .X(_04756_));
 sky130_fd_sc_hd__a211oi_1 _11941_ (.A1(_04652_),
    .A2(_04653_),
    .B1(_04755_),
    .C1(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__o211a_1 _11942_ (.A1(_04755_),
    .A2(_04756_),
    .B1(_04652_),
    .C1(_04653_),
    .X(_04758_));
 sky130_fd_sc_hd__o211a_1 _11943_ (.A1(_04757_),
    .A2(_04758_),
    .B1(_04604_),
    .C1(_04610_),
    .X(_04759_));
 sky130_fd_sc_hd__a211o_1 _11944_ (.A1(_04604_),
    .A2(_04610_),
    .B1(_04757_),
    .C1(_04758_),
    .X(_04760_));
 sky130_fd_sc_hd__nand2b_1 _11945_ (.A_N(_04759_),
    .B(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__o21ba_1 _11946_ (.A1(_04612_),
    .A2(_04613_),
    .B1_N(_04620_),
    .X(_04762_));
 sky130_fd_sc_hd__o21ai_1 _11947_ (.A1(_04761_),
    .A2(_04762_),
    .B1(_03133_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _11948_ (.A1(_04761_),
    .A2(_04762_),
    .B1(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__a211o_1 _11949_ (.A1(_03315_),
    .A2(_04641_),
    .B1(_04651_),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a31o_4 _11950_ (.A1(_02752_),
    .A2(_04637_),
    .A3(_04639_),
    .B1(_04765_),
    .X(net71));
 sky130_fd_sc_hd__o211ai_1 _11951_ (.A1(_04547_),
    .A2(_04549_),
    .B1(_04742_),
    .C1(_04743_),
    .Y(_04766_));
 sky130_fd_sc_hd__a22o_1 _11952_ (.A1(_02862_),
    .A2(_05906_),
    .B1(_05981_),
    .B2(_02808_),
    .X(_04768_));
 sky130_fd_sc_hd__nand4_2 _11953_ (.A(_02808_),
    .B(_02851_),
    .C(_05895_),
    .D(_05970_),
    .Y(_04769_));
 sky130_fd_sc_hd__or2b_1 _11954_ (.A(_04661_),
    .B_N(_04659_),
    .X(_04770_));
 sky130_fd_sc_hd__a32o_1 _11955_ (.A1(_06610_),
    .A2(_05831_),
    .A3(_04656_),
    .B1(_04655_),
    .B2(_05959_),
    .X(_04771_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_00058_),
    .B(_03449_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand4_1 _11957_ (.A(_02905_),
    .B(_02959_),
    .C(_05767_),
    .D(_05820_),
    .Y(_04773_));
 sky130_fd_sc_hd__a22o_1 _11958_ (.A1(_00216_),
    .A2(_03247_),
    .B1(_05820_),
    .B2(_00217_),
    .X(_04774_));
 sky130_fd_sc_hd__nand3b_1 _11959_ (.A_N(_04772_),
    .B(_04773_),
    .C(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__a21bo_1 _11960_ (.A1(_04774_),
    .A2(_04773_),
    .B1_N(_04772_),
    .X(_04776_));
 sky130_fd_sc_hd__nand3_1 _11961_ (.A(_04771_),
    .B(_04775_),
    .C(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__a21o_1 _11962_ (.A1(_04775_),
    .A2(_04776_),
    .B1(_04771_),
    .X(_04779_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(_04665_),
    .B(_04667_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21o_1 _11964_ (.A1(_04777_),
    .A2(_04779_),
    .B1(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__nand3_1 _11965_ (.A(_04780_),
    .B(_04777_),
    .C(_04779_),
    .Y(_04782_));
 sky130_fd_sc_hd__a21bo_1 _11966_ (.A1(_04670_),
    .A2(_04669_),
    .B1_N(_04668_),
    .X(_04783_));
 sky130_fd_sc_hd__nand3_1 _11967_ (.A(_04781_),
    .B(_04782_),
    .C(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__a21o_1 _11968_ (.A1(_04781_),
    .A2(_04782_),
    .B1(_04783_),
    .X(_04785_));
 sky130_fd_sc_hd__a22oi_2 _11969_ (.A1(_03282_),
    .A2(_05380_),
    .B1(_05445_),
    .B2(_00124_),
    .Y(_04786_));
 sky130_fd_sc_hd__and4_1 _11970_ (.A(_00299_),
    .B(_00231_),
    .C(_00530_),
    .D(_06666_),
    .X(_04787_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(net114),
    .B(_03047_),
    .Y(_04788_));
 sky130_fd_sc_hd__or3_1 _11972_ (.A(_04786_),
    .B(_04787_),
    .C(_04788_),
    .X(_04790_));
 sky130_fd_sc_hd__o21ai_1 _11973_ (.A1(_04786_),
    .A2(_04787_),
    .B1(_04788_),
    .Y(_04791_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(_04790_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__a22oi_2 _11975_ (.A1(_00462_),
    .A2(_05563_),
    .B1(_05638_),
    .B2(_00237_),
    .Y(_04793_));
 sky130_fd_sc_hd__and4_1 _11976_ (.A(net118),
    .B(net117),
    .C(_06461_),
    .D(_05627_),
    .X(_04794_));
 sky130_fd_sc_hd__nand2_1 _11977_ (.A(_03152_),
    .B(_00398_),
    .Y(_04795_));
 sky130_fd_sc_hd__or3_1 _11978_ (.A(_04793_),
    .B(_04794_),
    .C(_04795_),
    .X(_04796_));
 sky130_fd_sc_hd__o21ai_1 _11979_ (.A1(_04793_),
    .A2(_04794_),
    .B1(_04795_),
    .Y(_04797_));
 sky130_fd_sc_hd__o21bai_1 _11980_ (.A1(_04684_),
    .A2(_04686_),
    .B1_N(_04685_),
    .Y(_04798_));
 sky130_fd_sc_hd__and3_1 _11981_ (.A(_04796_),
    .B(_04797_),
    .C(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__a21oi_1 _11982_ (.A1(_04796_),
    .A2(_04797_),
    .B1(_04798_),
    .Y(_04801_));
 sky130_fd_sc_hd__nor2_1 _11983_ (.A(_04799_),
    .B(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__xnor2_2 _11984_ (.A(_04792_),
    .B(_04802_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21oi_1 _11985_ (.A1(_04784_),
    .A2(_04785_),
    .B1(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__and3_1 _11986_ (.A(_04803_),
    .B(_04784_),
    .C(_04785_),
    .X(_04805_));
 sky130_fd_sc_hd__nor3_1 _11987_ (.A(_04770_),
    .B(_04804_),
    .C(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__o21a_1 _11988_ (.A1(_04804_),
    .A2(_04805_),
    .B1(_04770_),
    .X(_04807_));
 sky130_fd_sc_hd__a211o_1 _11989_ (.A1(_04675_),
    .A2(_04695_),
    .B1(_04806_),
    .C1(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__o211ai_1 _11990_ (.A1(_04806_),
    .A2(_04807_),
    .B1(_04675_),
    .C1(_04695_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand4_2 _11991_ (.A(_04768_),
    .B(_04769_),
    .C(_04808_),
    .D(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__a22o_1 _11992_ (.A1(_04768_),
    .A2(_04769_),
    .B1(_04808_),
    .B2(_04809_),
    .X(_04812_));
 sky130_fd_sc_hd__and3_1 _11993_ (.A(_04700_),
    .B(_04810_),
    .C(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__a21oi_1 _11994_ (.A1(_04810_),
    .A2(_04812_),
    .B1(_04700_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_1 _11995_ (.A(_04740_),
    .B(_04742_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_1 _11996_ (.A(_04510_),
    .B(_04694_),
    .C(_04695_),
    .Y(_04816_));
 sky130_fd_sc_hd__and3_1 _11997_ (.A(net112),
    .B(_03593_),
    .C(_04961_),
    .X(_04817_));
 sky130_fd_sc_hd__a22o_1 _11998_ (.A1(_03593_),
    .A2(_04961_),
    .B1(_06584_),
    .B2(_03539_),
    .X(_04818_));
 sky130_fd_sc_hd__a21bo_1 _11999_ (.A1(_00421_),
    .A2(_04817_),
    .B1_N(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _12000_ (.A(_03658_),
    .B(_00550_),
    .Y(_04820_));
 sky130_fd_sc_hd__xor2_1 _12001_ (.A(_04819_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__a32o_1 _12002_ (.A1(_02965_),
    .A2(_04854_),
    .A3(_04708_),
    .B1(_04707_),
    .B2(_04983_),
    .X(_04822_));
 sky130_fd_sc_hd__xor2_1 _12003_ (.A(_04821_),
    .B(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__and2_1 _12004_ (.A(_03722_),
    .B(_04854_),
    .X(_04824_));
 sky130_fd_sc_hd__xnor2_1 _12005_ (.A(_04823_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__and2_1 _12006_ (.A(_04711_),
    .B(_04712_),
    .X(_04826_));
 sky130_fd_sc_hd__a21oi_1 _12007_ (.A1(_04713_),
    .A2(_04715_),
    .B1(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__xnor2_1 _12008_ (.A(_04825_),
    .B(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2_1 _12009_ (.A(net61),
    .B(_04800_),
    .Y(_04829_));
 sky130_fd_sc_hd__xor2_2 _12010_ (.A(_04828_),
    .B(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__a21o_1 _12011_ (.A1(_04683_),
    .A2(_04691_),
    .B1(_04690_),
    .X(_04831_));
 sky130_fd_sc_hd__and4_1 _12012_ (.A(_03217_),
    .B(_03271_),
    .C(_06562_),
    .D(_06476_),
    .X(_04833_));
 sky130_fd_sc_hd__a31o_1 _12013_ (.A1(_00270_),
    .A2(_06561_),
    .A3(_04679_),
    .B1(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__a22o_1 _12014_ (.A1(_03432_),
    .A2(_06517_),
    .B1(_06518_),
    .B2(_00278_),
    .X(_04835_));
 sky130_fd_sc_hd__nand4_2 _12015_ (.A(_03378_),
    .B(_00279_),
    .C(_05187_),
    .D(_05252_),
    .Y(_04836_));
 sky130_fd_sc_hd__a22o_1 _12016_ (.A1(_00292_),
    .A2(_00534_),
    .B1(_04835_),
    .B2(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__nand4_2 _12017_ (.A(_00283_),
    .B(_00423_),
    .C(_04835_),
    .D(_04836_),
    .Y(_04838_));
 sky130_fd_sc_hd__nand3_2 _12018_ (.A(_04834_),
    .B(_04837_),
    .C(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__a21o_1 _12019_ (.A1(_04837_),
    .A2(_04838_),
    .B1(_04834_),
    .X(_04840_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(_04727_),
    .B(_04729_),
    .Y(_04841_));
 sky130_fd_sc_hd__a21o_1 _12021_ (.A1(_04839_),
    .A2(_04840_),
    .B1(_04841_),
    .X(_04842_));
 sky130_fd_sc_hd__nand3_2 _12022_ (.A(_04841_),
    .B(_04839_),
    .C(_04840_),
    .Y(_04844_));
 sky130_fd_sc_hd__and3_1 _12023_ (.A(_04831_),
    .B(_04842_),
    .C(_04844_),
    .X(_04845_));
 sky130_fd_sc_hd__a21oi_1 _12024_ (.A1(_04842_),
    .A2(_04844_),
    .B1(_04831_),
    .Y(_04846_));
 sky130_fd_sc_hd__a211o_1 _12025_ (.A1(_04730_),
    .A2(_04734_),
    .B1(_04845_),
    .C1(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__o211ai_1 _12026_ (.A1(_04845_),
    .A2(_04846_),
    .B1(_04730_),
    .C1(_04734_),
    .Y(_04848_));
 sky130_fd_sc_hd__o211ai_2 _12027_ (.A1(_04735_),
    .A2(_04738_),
    .B1(_04847_),
    .C1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__a211o_1 _12028_ (.A1(_04847_),
    .A2(_04848_),
    .B1(_04735_),
    .C1(_04738_),
    .X(_04850_));
 sky130_fd_sc_hd__and3_1 _12029_ (.A(_04830_),
    .B(_04849_),
    .C(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__a21oi_1 _12030_ (.A1(_04849_),
    .A2(_04850_),
    .B1(_04830_),
    .Y(_04852_));
 sky130_fd_sc_hd__a211o_1 _12031_ (.A1(_04816_),
    .A2(_04698_),
    .B1(_04851_),
    .C1(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__o211ai_1 _12032_ (.A1(_04851_),
    .A2(_04852_),
    .B1(_04816_),
    .C1(_04698_),
    .Y(_04855_));
 sky130_fd_sc_hd__and3_1 _12033_ (.A(_04815_),
    .B(_04853_),
    .C(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__a21oi_1 _12034_ (.A1(_04853_),
    .A2(_04855_),
    .B1(_04815_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor4_2 _12035_ (.A(_04813_),
    .B(_04814_),
    .C(_04856_),
    .D(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__o22a_1 _12036_ (.A1(_04813_),
    .A2(_04814_),
    .B1(_04856_),
    .B2(_04857_),
    .X(_04859_));
 sky130_fd_sc_hd__a211oi_1 _12037_ (.A1(_04702_),
    .A2(_04749_),
    .B1(_04858_),
    .C1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__o211a_1 _12038_ (.A1(_04858_),
    .A2(_04859_),
    .B1(_04702_),
    .C1(_04749_),
    .X(_04861_));
 sky130_fd_sc_hd__a211o_2 _12039_ (.A1(_04766_),
    .A2(_04746_),
    .B1(_04860_),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__o211ai_2 _12040_ (.A1(_04860_),
    .A2(_04861_),
    .B1(_04766_),
    .C1(_04746_),
    .Y(_04863_));
 sky130_fd_sc_hd__o211ai_4 _12041_ (.A1(_04751_),
    .A2(_04753_),
    .B1(_04862_),
    .C1(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__a211o_2 _12042_ (.A1(_04862_),
    .A2(_04863_),
    .B1(_04751_),
    .C1(_04753_),
    .X(_04866_));
 sky130_fd_sc_hd__a31o_1 _12043_ (.A1(_03820_),
    .A2(_04736_),
    .A3(_04719_),
    .B1(_04717_),
    .X(_04867_));
 sky130_fd_sc_hd__nand3_1 _12044_ (.A(_04864_),
    .B(_04866_),
    .C(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__a21o_1 _12045_ (.A1(_04864_),
    .A2(_04866_),
    .B1(_04867_),
    .X(_04869_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(_04868_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_1 _12047_ (.A(_04755_),
    .B(_04757_),
    .Y(_04871_));
 sky130_fd_sc_hd__xnor2_1 _12048_ (.A(_04870_),
    .B(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__nor3_1 _12049_ (.A(_04614_),
    .B(_04615_),
    .C(_04761_),
    .Y(_04873_));
 sky130_fd_sc_hd__inv_2 _12050_ (.A(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__or3_1 _12051_ (.A(_04612_),
    .B(_04613_),
    .C(_04759_),
    .X(_04875_));
 sky130_fd_sc_hd__o311ai_1 _12052_ (.A1(_04614_),
    .A2(_04616_),
    .A3(_04761_),
    .B1(_04875_),
    .C1(_04760_),
    .Y(_04877_));
 sky130_fd_sc_hd__o21ba_1 _12053_ (.A1(_04322_),
    .A2(_04874_),
    .B1_N(_04877_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _12054_ (.A(_04872_),
    .B(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__or2_1 _12055_ (.A(_04872_),
    .B(_04878_),
    .X(_04880_));
 sky130_fd_sc_hd__and2_1 _12056_ (.A(_02575_),
    .B(_02579_),
    .X(_04881_));
 sky130_fd_sc_hd__o21ai_1 _12057_ (.A1(_02575_),
    .A2(_02579_),
    .B1(_03315_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21a_1 _12058_ (.A1(_02871_),
    .A2(_04647_),
    .B1(_01233_),
    .X(_04883_));
 sky130_fd_sc_hd__xnor2_1 _12059_ (.A(_02844_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__a211oi_1 _12060_ (.A1(_02705_),
    .A2(_00566_),
    .B1(_03306_),
    .C1(_02843_),
    .Y(_04885_));
 sky130_fd_sc_hd__a221o_1 _12061_ (.A1(_00566_),
    .A2(_02745_),
    .B1(_04642_),
    .B2(_04671_),
    .C1(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__a2bb2o_1 _12062_ (.A1_N(_04736_),
    .A2_N(_02727_),
    .B1(_02718_),
    .B2(_04800_),
    .X(_04887_));
 sky130_fd_sc_hd__a221o_1 _12063_ (.A1(\FuI.Integer[12] ),
    .A2(_02931_),
    .B1(_02938_),
    .B2(\AuI.result[12] ),
    .C1(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__a211o_1 _12064_ (.A1(\MuI.result[12] ),
    .A2(_02739_),
    .B1(_04886_),
    .C1(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__a21oi_1 _12065_ (.A1(_04161_),
    .A2(_04884_),
    .B1(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__o21ai_2 _12066_ (.A1(_04881_),
    .A2(_04882_),
    .B1(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21bai_1 _12067_ (.A1(_02869_),
    .A2(_04634_),
    .B1_N(_02870_),
    .Y(_04892_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(_04892_),
    .A1(_02893_),
    .S(_02926_),
    .X(_04893_));
 sky130_fd_sc_hd__a21oi_1 _12069_ (.A1(_02844_),
    .A2(_04893_),
    .B1(_02713_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21a_1 _12070_ (.A1(_02844_),
    .A2(_04893_),
    .B1(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__a311o_4 _12071_ (.A1(_03134_),
    .A2(_04879_),
    .A3(_04880_),
    .B1(_04891_),
    .C1(_04895_),
    .X(net72));
 sky130_fd_sc_hd__or2b_1 _12072_ (.A(_04736_),
    .B_N(_02765_),
    .X(_04897_));
 sky130_fd_sc_hd__o21a_1 _12073_ (.A1(_02844_),
    .A2(_04892_),
    .B1(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__clkinv_2 _12074_ (.A(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__mux2_1 _12075_ (.A0(_04899_),
    .A1(_02896_),
    .S(_02928_),
    .X(_04900_));
 sky130_fd_sc_hd__xnor2_1 _12076_ (.A(_02848_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__or2_1 _12077_ (.A(_04825_),
    .B(_04827_),
    .X(_04902_));
 sky130_fd_sc_hd__or2_1 _12078_ (.A(_04828_),
    .B(_04829_),
    .X(_04903_));
 sky130_fd_sc_hd__a211o_1 _12079_ (.A1(_04702_),
    .A2(_04749_),
    .B1(_04858_),
    .C1(_04859_),
    .X(_04904_));
 sky130_fd_sc_hd__inv_2 _12080_ (.A(_04856_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_02862_),
    .B(_05981_),
    .Y(_04906_));
 sky130_fd_sc_hd__a22oi_1 _12082_ (.A1(_00216_),
    .A2(_05820_),
    .B1(_03444_),
    .B2(_00217_),
    .Y(_04908_));
 sky130_fd_sc_hd__and4_1 _12083_ (.A(_02894_),
    .B(_00046_),
    .C(_00783_),
    .D(_05884_),
    .X(_04909_));
 sky130_fd_sc_hd__o2bb2a_1 _12084_ (.A1_N(_00444_),
    .A2_N(_05767_),
    .B1(_04908_),
    .B2(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__and4bb_1 _12085_ (.A_N(_04908_),
    .B_N(_04909_),
    .C(_00058_),
    .D(_05767_),
    .X(_04911_));
 sky130_fd_sc_hd__nor2_1 _12086_ (.A(_04910_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__xnor2_1 _12087_ (.A(_04769_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_1 _12088_ (.A(_04773_),
    .B(_04775_),
    .Y(_04914_));
 sky130_fd_sc_hd__xnor2_1 _12089_ (.A(_04913_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__and2_1 _12090_ (.A(_04777_),
    .B(_04782_),
    .X(_04916_));
 sky130_fd_sc_hd__xnor2_1 _12091_ (.A(_04915_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__a22oi_1 _12092_ (.A1(_00727_),
    .A2(_06546_),
    .B1(_03051_),
    .B2(_00728_),
    .Y(_04919_));
 sky130_fd_sc_hd__and4_1 _12093_ (.A(_03228_),
    .B(_03282_),
    .C(_05445_),
    .D(_05509_),
    .X(_04920_));
 sky130_fd_sc_hd__nor2_1 _12094_ (.A(_04919_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(_03324_),
    .B(_05391_),
    .Y(_04922_));
 sky130_fd_sc_hd__xnor2_1 _12096_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(_00262_),
    .B(_03071_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand4_1 _12098_ (.A(_00921_),
    .B(_01206_),
    .C(_05649_),
    .D(_03449_),
    .Y(_04925_));
 sky130_fd_sc_hd__a22o_1 _12099_ (.A1(_01206_),
    .A2(_03425_),
    .B1(_05702_),
    .B2(_00921_),
    .X(_04926_));
 sky130_fd_sc_hd__nand3b_1 _12100_ (.A_N(_04924_),
    .B(_04925_),
    .C(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__a21bo_1 _12101_ (.A1(_04926_),
    .A2(_04925_),
    .B1_N(_04924_),
    .X(_04928_));
 sky130_fd_sc_hd__o21bai_1 _12102_ (.A1(_04793_),
    .A2(_04795_),
    .B1_N(_04794_),
    .Y(_04930_));
 sky130_fd_sc_hd__and3_1 _12103_ (.A(_04927_),
    .B(_04928_),
    .C(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__a21o_1 _12104_ (.A1(_04927_),
    .A2(_04928_),
    .B1(_04930_),
    .X(_04932_));
 sky130_fd_sc_hd__and2b_1 _12105_ (.A_N(_04931_),
    .B(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__xnor2_1 _12106_ (.A(_04923_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__xor2_1 _12107_ (.A(_04917_),
    .B(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a21boi_1 _12108_ (.A1(_04803_),
    .A2(_04785_),
    .B1_N(_04784_),
    .Y(_04936_));
 sky130_fd_sc_hd__xnor2_1 _12109_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__xor2_1 _12110_ (.A(_04906_),
    .B(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__xor2_1 _12111_ (.A(_04810_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__inv_2 _12112_ (.A(_04851_),
    .Y(_04941_));
 sky130_fd_sc_hd__or3_1 _12113_ (.A(_04770_),
    .B(_04804_),
    .C(_04805_),
    .X(_04942_));
 sky130_fd_sc_hd__and3_1 _12114_ (.A(net112),
    .B(_03593_),
    .C(_05025_),
    .X(_04943_));
 sky130_fd_sc_hd__a22o_1 _12115_ (.A1(_03593_),
    .A2(_05025_),
    .B1(_06623_),
    .B2(net112),
    .X(_04944_));
 sky130_fd_sc_hd__a21bo_1 _12116_ (.A1(_00534_),
    .A2(_04943_),
    .B1_N(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__nand2_1 _12117_ (.A(_06439_),
    .B(_00197_),
    .Y(_04946_));
 sky130_fd_sc_hd__xor2_1 _12118_ (.A(_04945_),
    .B(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__a32o_1 _12119_ (.A1(_03658_),
    .A2(_04918_),
    .A3(_04818_),
    .B1(_04817_),
    .B2(_05047_),
    .X(_04948_));
 sky130_fd_sc_hd__xor2_2 _12120_ (.A(_04947_),
    .B(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__and2_1 _12121_ (.A(net60),
    .B(_04918_),
    .X(_04950_));
 sky130_fd_sc_hd__xnor2_2 _12122_ (.A(_04949_),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__and2_1 _12123_ (.A(_04821_),
    .B(_04822_),
    .X(_04952_));
 sky130_fd_sc_hd__a21oi_2 _12124_ (.A1(_04823_),
    .A2(_04824_),
    .B1(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__xor2_2 _12125_ (.A(_04951_),
    .B(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__nand2_1 _12126_ (.A(net61),
    .B(_04854_),
    .Y(_04955_));
 sky130_fd_sc_hd__xnor2_2 _12127_ (.A(_04954_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand3_1 _12128_ (.A(_04831_),
    .B(_04842_),
    .C(_04844_),
    .Y(_04957_));
 sky130_fd_sc_hd__o21bai_1 _12129_ (.A1(_04792_),
    .A2(_04801_),
    .B1_N(_04799_),
    .Y(_04958_));
 sky130_fd_sc_hd__o21bai_1 _12130_ (.A1(_04786_),
    .A2(_04788_),
    .B1_N(_04787_),
    .Y(_04959_));
 sky130_fd_sc_hd__a22o_1 _12131_ (.A1(_00279_),
    .A2(_05252_),
    .B1(_00412_),
    .B2(_00278_),
    .X(_04960_));
 sky130_fd_sc_hd__nand4_2 _12132_ (.A(_03378_),
    .B(_00289_),
    .C(_05252_),
    .D(_05316_),
    .Y(_04962_));
 sky130_fd_sc_hd__a22o_1 _12133_ (.A1(_00292_),
    .A2(_00002_),
    .B1(_04960_),
    .B2(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__nand4_2 _12134_ (.A(_00283_),
    .B(_05198_),
    .C(_04960_),
    .D(_04962_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand3_1 _12135_ (.A(_04959_),
    .B(_04963_),
    .C(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__a21o_1 _12136_ (.A1(_04963_),
    .A2(_04964_),
    .B1(_04959_),
    .X(_04966_));
 sky130_fd_sc_hd__nand2_1 _12137_ (.A(_04836_),
    .B(_04838_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21o_1 _12138_ (.A1(_04965_),
    .A2(_04966_),
    .B1(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__nand3_1 _12139_ (.A(_04967_),
    .B(_04965_),
    .C(_04966_),
    .Y(_04969_));
 sky130_fd_sc_hd__and3_1 _12140_ (.A(_04958_),
    .B(_04968_),
    .C(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__a21oi_1 _12141_ (.A1(_04968_),
    .A2(_04969_),
    .B1(_04958_),
    .Y(_04971_));
 sky130_fd_sc_hd__a211oi_2 _12142_ (.A1(_04839_),
    .A2(_04844_),
    .B1(_04970_),
    .C1(_04971_),
    .Y(_04973_));
 sky130_fd_sc_hd__o211a_1 _12143_ (.A1(_04970_),
    .A2(_04971_),
    .B1(_04839_),
    .C1(_04844_),
    .X(_04974_));
 sky130_fd_sc_hd__a211o_1 _12144_ (.A1(_04957_),
    .A2(_04847_),
    .B1(_04973_),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o211ai_1 _12145_ (.A1(_04973_),
    .A2(_04974_),
    .B1(_04957_),
    .C1(_04847_),
    .Y(_04976_));
 sky130_fd_sc_hd__and3_1 _12146_ (.A(_04956_),
    .B(_04975_),
    .C(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__a21oi_1 _12147_ (.A1(_04975_),
    .A2(_04976_),
    .B1(_04956_),
    .Y(_04978_));
 sky130_fd_sc_hd__a211oi_1 _12148_ (.A1(_04942_),
    .A2(_04808_),
    .B1(_04977_),
    .C1(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__o211a_1 _12149_ (.A1(_04977_),
    .A2(_04978_),
    .B1(_04942_),
    .C1(_04808_),
    .X(_04980_));
 sky130_fd_sc_hd__a211o_2 _12150_ (.A1(_04849_),
    .A2(_04941_),
    .B1(_04979_),
    .C1(_04980_),
    .X(_04981_));
 sky130_fd_sc_hd__o211ai_1 _12151_ (.A1(_04979_),
    .A2(_04980_),
    .B1(_04849_),
    .C1(_04941_),
    .Y(_04982_));
 sky130_fd_sc_hd__and3_1 _12152_ (.A(_04939_),
    .B(_04981_),
    .C(_04982_),
    .X(_04984_));
 sky130_fd_sc_hd__a21oi_1 _12153_ (.A1(_04981_),
    .A2(_04982_),
    .B1(_04939_),
    .Y(_04985_));
 sky130_fd_sc_hd__nor2_1 _12154_ (.A(_04984_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21a_2 _12155_ (.A1(_04813_),
    .A2(_04858_),
    .B1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__nor3_2 _12156_ (.A(_04813_),
    .B(_04858_),
    .C(_04986_),
    .Y(_04988_));
 sky130_fd_sc_hd__a211oi_4 _12157_ (.A1(_04853_),
    .A2(_04905_),
    .B1(_04987_),
    .C1(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__o211a_1 _12158_ (.A1(_04987_),
    .A2(_04988_),
    .B1(_04853_),
    .C1(_04905_),
    .X(_04990_));
 sky130_fd_sc_hd__a211oi_4 _12159_ (.A1(_04904_),
    .A2(_04862_),
    .B1(_04989_),
    .C1(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__o211a_2 _12160_ (.A1(_04989_),
    .A2(_04990_),
    .B1(_04904_),
    .C1(_04862_),
    .X(_04992_));
 sky130_fd_sc_hd__a211oi_2 _12161_ (.A1(_04902_),
    .A2(_04903_),
    .B1(_04991_),
    .C1(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__o211a_1 _12162_ (.A1(_04991_),
    .A2(_04992_),
    .B1(_04902_),
    .C1(_04903_),
    .X(_04995_));
 sky130_fd_sc_hd__a211oi_1 _12163_ (.A1(_04864_),
    .A2(_04868_),
    .B1(_04993_),
    .C1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__o211a_1 _12164_ (.A1(_04993_),
    .A2(_04995_),
    .B1(_04864_),
    .C1(_04868_),
    .X(_04997_));
 sky130_fd_sc_hd__or2_1 _12165_ (.A(_04996_),
    .B(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__nor2_1 _12166_ (.A(_04870_),
    .B(_04871_),
    .Y(_04999_));
 sky130_fd_sc_hd__and2b_1 _12167_ (.A_N(_04999_),
    .B(_04880_),
    .X(_05000_));
 sky130_fd_sc_hd__o21ai_1 _12168_ (.A1(_04998_),
    .A2(_05000_),
    .B1(_03134_),
    .Y(_05001_));
 sky130_fd_sc_hd__a21oi_1 _12169_ (.A1(_04998_),
    .A2(_05000_),
    .B1(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21bai_1 _12170_ (.A1(_02843_),
    .A2(_04883_),
    .B1_N(_00566_),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _12171_ (.A(_02848_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__o21a_1 _12172_ (.A1(_02848_),
    .A2(_05003_),
    .B1(_04161_),
    .X(_05006_));
 sky130_fd_sc_hd__o21ai_1 _12173_ (.A1(_02581_),
    .A2(_04881_),
    .B1(_02447_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _12174_ (.A(_02444_),
    .B(_02446_),
    .Y(_05008_));
 sky130_fd_sc_hd__a211o_1 _12175_ (.A1(_02447_),
    .A2(_05008_),
    .B1(_02581_),
    .C1(_04881_),
    .X(_05009_));
 sky130_fd_sc_hd__a2bb2o_1 _12176_ (.A1_N(_04800_),
    .A2_N(_02941_),
    .B1(_02938_),
    .B2(\AuI.result[13] ),
    .X(_05010_));
 sky130_fd_sc_hd__a22o_1 _12177_ (.A1(\MuI.result[13] ),
    .A2(_02736_),
    .B1(_02944_),
    .B2(_04736_),
    .X(_05011_));
 sky130_fd_sc_hd__a221o_1 _12178_ (.A1(_00555_),
    .A2(_02743_),
    .B1(_02848_),
    .B2(_04011_),
    .C1(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__a221o_1 _12179_ (.A1(\FuI.Integer[13] ),
    .A2(_02931_),
    .B1(_03675_),
    .B2(_04865_),
    .C1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a211o_1 _12180_ (.A1(_02808_),
    .A2(_02724_),
    .B1(_05010_),
    .C1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__a31o_1 _12181_ (.A1(_05007_),
    .A2(_03314_),
    .A3(_05009_),
    .B1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__a21o_1 _12182_ (.A1(_05004_),
    .A2(_05006_),
    .B1(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__a211o_4 _12183_ (.A1(_02751_),
    .A2(_04901_),
    .B1(_05002_),
    .C1(_05016_),
    .X(net73));
 sky130_fd_sc_hd__a21o_1 _12184_ (.A1(_02845_),
    .A2(_04898_),
    .B1(_02846_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(_05017_),
    .A1(_02897_),
    .S(_02928_),
    .X(_05018_));
 sky130_fd_sc_hd__or2_1 _12186_ (.A(_02795_),
    .B(_05018_),
    .X(_05019_));
 sky130_fd_sc_hd__nand2_1 _12187_ (.A(_02795_),
    .B(_05018_),
    .Y(_05020_));
 sky130_fd_sc_hd__and3_1 _12188_ (.A(_02402_),
    .B(_05008_),
    .C(_05007_),
    .X(_05021_));
 sky130_fd_sc_hd__o21a_1 _12189_ (.A1(_02862_),
    .A2(_04865_),
    .B1(_02722_),
    .X(_05022_));
 sky130_fd_sc_hd__a32o_1 _12190_ (.A1(_02862_),
    .A2(_04865_),
    .A3(_02745_),
    .B1(_02719_),
    .B2(_04929_),
    .X(_05023_));
 sky130_fd_sc_hd__a211o_1 _12191_ (.A1(_04800_),
    .A2(_04642_),
    .B1(_05022_),
    .C1(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__a2bb2o_1 _12192_ (.A1_N(_04865_),
    .A2_N(_02728_),
    .B1(_02931_),
    .B2(\FuI.Integer[14] ),
    .X(_05026_));
 sky130_fd_sc_hd__a221o_1 _12193_ (.A1(\MuI.result[14] ),
    .A2(_02739_),
    .B1(_03494_),
    .B2(_02795_),
    .C1(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__a21o_1 _12194_ (.A1(_02848_),
    .A2(_05003_),
    .B1(_00555_),
    .X(_05028_));
 sky130_fd_sc_hd__nand2_1 _12195_ (.A(_02795_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__or2_1 _12196_ (.A(_02795_),
    .B(_05028_),
    .X(_05030_));
 sky130_fd_sc_hd__a32o_1 _12197_ (.A1(_02935_),
    .A2(_05029_),
    .A3(_05030_),
    .B1(_02732_),
    .B2(\AuI.result[14] ),
    .X(_05031_));
 sky130_fd_sc_hd__nor3_1 _12198_ (.A(_05024_),
    .B(_05027_),
    .C(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nor2_1 _12199_ (.A(_04951_),
    .B(_04953_),
    .Y(_05033_));
 sky130_fd_sc_hd__and3_1 _12200_ (.A(_03820_),
    .B(_04865_),
    .C(_04954_),
    .X(_05034_));
 sky130_fd_sc_hd__a211o_1 _12201_ (.A1(_04942_),
    .A2(_04808_),
    .B1(_04977_),
    .C1(_04978_),
    .X(_05035_));
 sky130_fd_sc_hd__nor2_1 _12202_ (.A(_04810_),
    .B(_04938_),
    .Y(_05037_));
 sky130_fd_sc_hd__or2b_1 _12203_ (.A(_04906_),
    .B_N(_04937_),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(_02959_),
    .B(_03444_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(_02905_),
    .B(_05959_),
    .Y(_05040_));
 sky130_fd_sc_hd__and2_1 _12206_ (.A(_00029_),
    .B(_00153_),
    .X(_05041_));
 sky130_fd_sc_hd__and3_1 _12207_ (.A(_00217_),
    .B(_05948_),
    .C(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a21oi_1 _12208_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _12209_ (.A(_03024_),
    .B(_05831_),
    .Y(_05044_));
 sky130_fd_sc_hd__xnor2_1 _12210_ (.A(_05043_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nor2_1 _12211_ (.A(_04909_),
    .B(_04911_),
    .Y(_05046_));
 sky130_fd_sc_hd__xnor2_1 _12212_ (.A(_05045_),
    .B(_05046_),
    .Y(_05048_));
 sky130_fd_sc_hd__and2b_1 _12213_ (.A_N(_04769_),
    .B(_04912_),
    .X(_05049_));
 sky130_fd_sc_hd__a21oi_1 _12214_ (.A1(_04913_),
    .A2(_04914_),
    .B1(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__xnor2_1 _12215_ (.A(_05048_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_2 _12216_ (.A(_03335_),
    .B(_05456_),
    .Y(_05052_));
 sky130_fd_sc_hd__a22oi_1 _12217_ (.A1(_00727_),
    .A2(_03051_),
    .B1(_03071_),
    .B2(_00728_),
    .Y(_05053_));
 sky130_fd_sc_hd__and4_1 _12218_ (.A(_03228_),
    .B(_03282_),
    .C(_05509_),
    .D(_05574_),
    .X(_05054_));
 sky130_fd_sc_hd__nor2_1 _12219_ (.A(_05053_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_1 _12220_ (.A(_05052_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _12221_ (.A(_03163_),
    .B(_03425_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand4_1 _12222_ (.A(_00921_),
    .B(_00132_),
    .C(_05702_),
    .D(_03247_),
    .Y(_05059_));
 sky130_fd_sc_hd__a22o_1 _12223_ (.A1(_00132_),
    .A2(_00163_),
    .B1(_00385_),
    .B2(_00133_),
    .X(_05060_));
 sky130_fd_sc_hd__nand3b_1 _12224_ (.A_N(_05057_),
    .B(_05059_),
    .C(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__a21bo_1 _12225_ (.A1(_05060_),
    .A2(_05059_),
    .B1_N(_05057_),
    .X(_05062_));
 sky130_fd_sc_hd__nand2_1 _12226_ (.A(_05061_),
    .B(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _12227_ (.A(_04925_),
    .B(_04927_),
    .Y(_05064_));
 sky130_fd_sc_hd__xnor2_1 _12228_ (.A(_05063_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__xnor2_1 _12229_ (.A(_05056_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_2 _12230_ (.A(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _12231_ (.A(_05051_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__or2_1 _12232_ (.A(_05051_),
    .B(_05067_),
    .X(_05070_));
 sky130_fd_sc_hd__nand2_1 _12233_ (.A(_05068_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__or2_1 _12234_ (.A(_04915_),
    .B(_04916_),
    .X(_05072_));
 sky130_fd_sc_hd__o21ai_1 _12235_ (.A1(_04917_),
    .A2(_04934_),
    .B1(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__xor2_1 _12236_ (.A(_05071_),
    .B(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__xor2_1 _12237_ (.A(_05038_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__inv_2 _12238_ (.A(_04977_),
    .Y(_05076_));
 sky130_fd_sc_hd__or2b_1 _12239_ (.A(_04936_),
    .B_N(_04935_),
    .X(_05077_));
 sky130_fd_sc_hd__a22oi_2 _12240_ (.A1(_06442_),
    .A2(_00423_),
    .B1(_00002_),
    .B2(_03550_),
    .Y(_05078_));
 sky130_fd_sc_hd__and4_1 _12241_ (.A(_06444_),
    .B(_06442_),
    .C(_00534_),
    .D(_06525_),
    .X(_05079_));
 sky130_fd_sc_hd__nor2_2 _12242_ (.A(_05078_),
    .B(_05079_),
    .Y(_05081_));
 sky130_fd_sc_hd__nand2_2 _12243_ (.A(_03658_),
    .B(_05047_),
    .Y(_05082_));
 sky130_fd_sc_hd__xnor2_4 _12244_ (.A(_05081_),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__a32o_2 _12245_ (.A1(_03525_),
    .A2(_04983_),
    .A3(_04944_),
    .B1(_04943_),
    .B2(_05123_),
    .X(_05084_));
 sky130_fd_sc_hd__xor2_4 _12246_ (.A(_05083_),
    .B(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__nand2_1 _12247_ (.A(_06429_),
    .B(_04983_),
    .Y(_05086_));
 sky130_fd_sc_hd__xor2_4 _12248_ (.A(_05085_),
    .B(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__and2_1 _12249_ (.A(_04947_),
    .B(_04948_),
    .X(_05088_));
 sky130_fd_sc_hd__a21oi_2 _12250_ (.A1(_04949_),
    .A2(_04950_),
    .B1(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__xnor2_4 _12251_ (.A(_05087_),
    .B(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_2 _12252_ (.A(_00502_),
    .B(_04918_),
    .Y(_05091_));
 sky130_fd_sc_hd__xor2_4 _12253_ (.A(_05090_),
    .B(_05091_),
    .X(_05092_));
 sky130_fd_sc_hd__a21o_1 _12254_ (.A1(_04923_),
    .A2(_04932_),
    .B1(_04931_),
    .X(_05093_));
 sky130_fd_sc_hd__o21bai_1 _12255_ (.A1(_04919_),
    .A2(_04922_),
    .B1_N(_04920_),
    .Y(_05094_));
 sky130_fd_sc_hd__a22o_1 _12256_ (.A1(_02980_),
    .A2(_03047_),
    .B1(_06477_),
    .B2(_00281_),
    .X(_05095_));
 sky130_fd_sc_hd__nand4_1 _12257_ (.A(_02983_),
    .B(_02984_),
    .C(_03047_),
    .D(_06477_),
    .Y(_05096_));
 sky130_fd_sc_hd__a22o_1 _12258_ (.A1(_03486_),
    .A2(_05262_),
    .B1(_05095_),
    .B2(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__nand4_1 _12259_ (.A(_02987_),
    .B(_05262_),
    .C(_05095_),
    .D(_05096_),
    .Y(_05098_));
 sky130_fd_sc_hd__nand3_2 _12260_ (.A(_05094_),
    .B(_05097_),
    .C(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__a21o_1 _12261_ (.A1(_05097_),
    .A2(_05098_),
    .B1(_05094_),
    .X(_05100_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_04962_),
    .B(_04964_),
    .Y(_05102_));
 sky130_fd_sc_hd__a21o_1 _12263_ (.A1(_05099_),
    .A2(_05100_),
    .B1(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__nand3_2 _12264_ (.A(_05102_),
    .B(_05099_),
    .C(_05100_),
    .Y(_05104_));
 sky130_fd_sc_hd__and3_1 _12265_ (.A(_05093_),
    .B(_05103_),
    .C(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__a21oi_1 _12266_ (.A1(_05103_),
    .A2(_05104_),
    .B1(_05093_),
    .Y(_05106_));
 sky130_fd_sc_hd__a211o_2 _12267_ (.A1(_04965_),
    .A2(_04969_),
    .B1(_05105_),
    .C1(_05106_),
    .X(_05107_));
 sky130_fd_sc_hd__o211ai_1 _12268_ (.A1(_05105_),
    .A2(_05106_),
    .B1(_04965_),
    .C1(_04969_),
    .Y(_05108_));
 sky130_fd_sc_hd__o211ai_2 _12269_ (.A1(_04970_),
    .A2(_04973_),
    .B1(_05107_),
    .C1(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__a211o_1 _12270_ (.A1(_05107_),
    .A2(_05108_),
    .B1(_04970_),
    .C1(_04973_),
    .X(_05110_));
 sky130_fd_sc_hd__and3_1 _12271_ (.A(_05092_),
    .B(_05109_),
    .C(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21oi_2 _12272_ (.A1(_05109_),
    .A2(_05110_),
    .B1(_05092_),
    .Y(_05113_));
 sky130_fd_sc_hd__nor3_4 _12273_ (.A(_05077_),
    .B(_05111_),
    .C(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__o21a_1 _12274_ (.A1(_05111_),
    .A2(_05113_),
    .B1(_05077_),
    .X(_05115_));
 sky130_fd_sc_hd__a211o_1 _12275_ (.A1(_04975_),
    .A2(_05076_),
    .B1(_05114_),
    .C1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o211ai_1 _12276_ (.A1(_05114_),
    .A2(_05115_),
    .B1(_04975_),
    .C1(_05076_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand3_1 _12277_ (.A(_05075_),
    .B(_05116_),
    .C(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__a21o_1 _12278_ (.A1(_05116_),
    .A2(_05117_),
    .B1(_05075_),
    .X(_05119_));
 sky130_fd_sc_hd__o211a_2 _12279_ (.A1(_05037_),
    .A2(_04984_),
    .B1(_05118_),
    .C1(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__a211oi_4 _12280_ (.A1(_05118_),
    .A2(_05119_),
    .B1(_05037_),
    .C1(_04984_),
    .Y(_05121_));
 sky130_fd_sc_hd__a211oi_4 _12281_ (.A1(_05035_),
    .A2(_04981_),
    .B1(_05120_),
    .C1(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__inv_2 _12282_ (.A(_05122_),
    .Y(_05124_));
 sky130_fd_sc_hd__o211ai_2 _12283_ (.A1(_05120_),
    .A2(_05121_),
    .B1(_05035_),
    .C1(_04981_),
    .Y(_05125_));
 sky130_fd_sc_hd__o211ai_4 _12284_ (.A1(_04987_),
    .A2(_04989_),
    .B1(_05124_),
    .C1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__a211o_2 _12285_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_04987_),
    .C1(_04989_),
    .X(_05127_));
 sky130_fd_sc_hd__o211ai_2 _12286_ (.A1(_05033_),
    .A2(_05034_),
    .B1(_05126_),
    .C1(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__a211o_1 _12287_ (.A1(_05126_),
    .A2(_05127_),
    .B1(_05033_),
    .C1(_05034_),
    .X(_05129_));
 sky130_fd_sc_hd__nand2_1 _12288_ (.A(_05128_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__nor2_1 _12289_ (.A(_04991_),
    .B(_04993_),
    .Y(_05131_));
 sky130_fd_sc_hd__xnor2_1 _12290_ (.A(_05130_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nor2_1 _12291_ (.A(_04999_),
    .B(_04996_),
    .Y(_05133_));
 sky130_fd_sc_hd__o32a_1 _12292_ (.A1(_04872_),
    .A2(_04878_),
    .A3(_04998_),
    .B1(_05133_),
    .B2(_04997_),
    .X(_05135_));
 sky130_fd_sc_hd__nor2_1 _12293_ (.A(_05132_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__nand2_1 _12294_ (.A(_05132_),
    .B(_05135_),
    .Y(_05137_));
 sky130_fd_sc_hd__or3b_1 _12295_ (.A(_05136_),
    .B(_06427_),
    .C_N(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__o311ai_2 _12296_ (.A1(_02584_),
    .A2(_04159_),
    .A3(_05021_),
    .B1(_05032_),
    .C1(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__a31o_2 _12297_ (.A1(_02752_),
    .A2(_05019_),
    .A3(_05020_),
    .B1(_05139_),
    .X(net74));
 sky130_fd_sc_hd__o21bai_1 _12298_ (.A1(_02795_),
    .A2(_05017_),
    .B1_N(_02792_),
    .Y(_05140_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(_05140_),
    .A1(_02898_),
    .S(_04635_),
    .X(_05141_));
 sky130_fd_sc_hd__nand2_1 _12300_ (.A(_02800_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__or2_1 _12301_ (.A(_02800_),
    .B(_05141_),
    .X(_05143_));
 sky130_fd_sc_hd__a211oi_2 _12302_ (.A1(_04975_),
    .A2(_05076_),
    .B1(_05114_),
    .C1(_05115_),
    .Y(_05145_));
 sky130_fd_sc_hd__nor2_1 _12303_ (.A(_05038_),
    .B(_05074_),
    .Y(_05146_));
 sky130_fd_sc_hd__and3_1 _12304_ (.A(_05075_),
    .B(_05116_),
    .C(_05117_),
    .X(_05147_));
 sky130_fd_sc_hd__or2b_1 _12305_ (.A(_05050_),
    .B_N(_05048_),
    .X(_05148_));
 sky130_fd_sc_hd__and2b_1 _12306_ (.A_N(_05046_),
    .B(_05045_),
    .X(_05149_));
 sky130_fd_sc_hd__and3_1 _12307_ (.A(_03013_),
    .B(_05831_),
    .C(_05043_),
    .X(_05150_));
 sky130_fd_sc_hd__nand2_1 _12308_ (.A(_03013_),
    .B(_05959_),
    .Y(_05151_));
 sky130_fd_sc_hd__a22o_1 _12309_ (.A1(_03013_),
    .A2(_05895_),
    .B1(_05959_),
    .B2(_02970_),
    .X(_05152_));
 sky130_fd_sc_hd__o21a_1 _12310_ (.A1(_05039_),
    .A2(_05151_),
    .B1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__o21ai_1 _12311_ (.A1(_05042_),
    .A2(_05150_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__or3_1 _12312_ (.A(_05042_),
    .B(_05150_),
    .C(_05153_),
    .X(_05156_));
 sky130_fd_sc_hd__and2_1 _12313_ (.A(_05154_),
    .B(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__xnor2_1 _12314_ (.A(_05149_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__a22oi_1 _12315_ (.A1(_00231_),
    .A2(_03424_),
    .B1(_00382_),
    .B2(_00299_),
    .Y(_05159_));
 sky130_fd_sc_hd__and4_1 _12316_ (.A(_03217_),
    .B(_03271_),
    .C(_05563_),
    .D(_05627_),
    .X(_05160_));
 sky130_fd_sc_hd__nor2_1 _12317_ (.A(_05159_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_1 _12318_ (.A(_03335_),
    .B(_05520_),
    .Y(_05162_));
 sky130_fd_sc_hd__xnor2_1 _12319_ (.A(_05161_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__a22oi_1 _12320_ (.A1(_00081_),
    .A2(_05756_),
    .B1(_00783_),
    .B2(_03056_),
    .Y(_05164_));
 sky130_fd_sc_hd__and4_1 _12321_ (.A(_00237_),
    .B(_00096_),
    .C(_05756_),
    .D(_00785_),
    .X(_05165_));
 sky130_fd_sc_hd__nor2_1 _12322_ (.A(_05164_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _12323_ (.A(_03163_),
    .B(_03449_),
    .Y(_05167_));
 sky130_fd_sc_hd__xnor2_2 _12324_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _12325_ (.A(_05059_),
    .B(_05061_),
    .Y(_05169_));
 sky130_fd_sc_hd__xor2_1 _12326_ (.A(_05168_),
    .B(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__and2_1 _12327_ (.A(_05163_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_1 _12328_ (.A(_05163_),
    .B(_05170_),
    .Y(_05172_));
 sky130_fd_sc_hd__or2_1 _12329_ (.A(_05171_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__nor2_1 _12330_ (.A(_05158_),
    .B(_05173_),
    .Y(_05174_));
 sky130_fd_sc_hd__and2_1 _12331_ (.A(_05158_),
    .B(_05173_),
    .X(_05175_));
 sky130_fd_sc_hd__or2_1 _12332_ (.A(_05174_),
    .B(_05175_),
    .X(_05177_));
 sky130_fd_sc_hd__a21o_1 _12333_ (.A1(_05148_),
    .A2(_05068_),
    .B1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__nand3_1 _12334_ (.A(_05148_),
    .B(_05068_),
    .C(_05177_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _12335_ (.A(_05178_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__a21boi_2 _12336_ (.A1(_05092_),
    .A2(_05110_),
    .B1_N(_05109_),
    .Y(_05181_));
 sky130_fd_sc_hd__or2b_1 _12337_ (.A(_05071_),
    .B_N(_05073_),
    .X(_05182_));
 sky130_fd_sc_hd__nand3_1 _12338_ (.A(_05093_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05183_));
 sky130_fd_sc_hd__a32o_1 _12339_ (.A1(_05061_),
    .A2(_05062_),
    .A3(_05064_),
    .B1(_05065_),
    .B2(_05056_),
    .X(_05184_));
 sky130_fd_sc_hd__a31o_1 _12340_ (.A1(_03335_),
    .A2(_05456_),
    .A3(_05055_),
    .B1(_05054_),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_1 _12341_ (.A1(_02984_),
    .A2(_06477_),
    .B1(_06546_),
    .B2(_03389_),
    .X(_05186_));
 sky130_fd_sc_hd__nand4_1 _12342_ (.A(_03389_),
    .B(_03454_),
    .C(_05391_),
    .D(_06546_),
    .Y(_05188_));
 sky130_fd_sc_hd__a22o_1 _12343_ (.A1(_03497_),
    .A2(_05327_),
    .B1(_05186_),
    .B2(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__nand4_1 _12344_ (.A(_03497_),
    .B(_05327_),
    .C(_05186_),
    .D(_05188_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand3_2 _12345_ (.A(_05185_),
    .B(_05189_),
    .C(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a21o_1 _12346_ (.A1(_05189_),
    .A2(_05190_),
    .B1(_05185_),
    .X(_05192_));
 sky130_fd_sc_hd__nand2_1 _12347_ (.A(_05096_),
    .B(_05098_),
    .Y(_05193_));
 sky130_fd_sc_hd__a21o_1 _12348_ (.A1(_05191_),
    .A2(_05192_),
    .B1(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__nand3_2 _12349_ (.A(_05193_),
    .B(_05191_),
    .C(_05192_),
    .Y(_05195_));
 sky130_fd_sc_hd__and3_2 _12350_ (.A(_05184_),
    .B(_05194_),
    .C(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__a21oi_2 _12351_ (.A1(_05194_),
    .A2(_05195_),
    .B1(_05184_),
    .Y(_05197_));
 sky130_fd_sc_hd__a211oi_4 _12352_ (.A1(_05099_),
    .A2(_05104_),
    .B1(_05196_),
    .C1(_05197_),
    .Y(_05199_));
 sky130_fd_sc_hd__o211a_1 _12353_ (.A1(_05196_),
    .A2(_05197_),
    .B1(_05099_),
    .C1(_05104_),
    .X(_05200_));
 sky130_fd_sc_hd__a211oi_4 _12354_ (.A1(_05183_),
    .A2(_05107_),
    .B1(_05199_),
    .C1(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hd__o211a_1 _12355_ (.A1(_05199_),
    .A2(_05200_),
    .B1(_05183_),
    .C1(_05107_),
    .X(_05202_));
 sky130_fd_sc_hd__a22oi_1 _12356_ (.A1(_06442_),
    .A2(_00002_),
    .B1(_06561_),
    .B2(_06444_),
    .Y(_05203_));
 sky130_fd_sc_hd__and4_1 _12357_ (.A(_00506_),
    .B(_00676_),
    .C(_06525_),
    .D(_06568_),
    .X(_05204_));
 sky130_fd_sc_hd__nor2_1 _12358_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(_06439_),
    .B(_05123_),
    .Y(_05206_));
 sky130_fd_sc_hd__xnor2_1 _12360_ (.A(_05205_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__o21ba_1 _12361_ (.A1(_05078_),
    .A2(_05082_),
    .B1_N(_05079_),
    .X(_05208_));
 sky130_fd_sc_hd__xnor2_1 _12362_ (.A(_05207_),
    .B(_05208_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand3_1 _12363_ (.A(_03733_),
    .B(_05047_),
    .C(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__a21o_1 _12364_ (.A1(_03733_),
    .A2(_05047_),
    .B1(_05210_),
    .X(_05212_));
 sky130_fd_sc_hd__nand2_1 _12365_ (.A(_05211_),
    .B(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__and2_1 _12366_ (.A(_05083_),
    .B(_05084_),
    .X(_05214_));
 sky130_fd_sc_hd__a31o_1 _12367_ (.A1(_03744_),
    .A2(_04983_),
    .A3(_05085_),
    .B1(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__xnor2_2 _12368_ (.A(_05213_),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _12369_ (.A(_03798_),
    .B(_04983_),
    .Y(_05217_));
 sky130_fd_sc_hd__xnor2_2 _12370_ (.A(_05216_),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nor3b_4 _12371_ (.A(_05201_),
    .B(_05202_),
    .C_N(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__o21ba_1 _12372_ (.A1(_05201_),
    .A2(_05202_),
    .B1_N(_05218_),
    .X(_05221_));
 sky130_fd_sc_hd__nor3_4 _12373_ (.A(_05182_),
    .B(_05219_),
    .C(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__o21a_1 _12374_ (.A1(_05219_),
    .A2(_05221_),
    .B1(_05182_),
    .X(_05223_));
 sky130_fd_sc_hd__nor3_4 _12375_ (.A(_05181_),
    .B(_05222_),
    .C(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__o21a_1 _12376_ (.A1(_05222_),
    .A2(_05223_),
    .B1(_05181_),
    .X(_05225_));
 sky130_fd_sc_hd__or3_2 _12377_ (.A(_05180_),
    .B(_05224_),
    .C(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__o21ai_2 _12378_ (.A1(_05224_),
    .A2(_05225_),
    .B1(_05180_),
    .Y(_05227_));
 sky130_fd_sc_hd__o211ai_4 _12379_ (.A1(_05146_),
    .A2(_05147_),
    .B1(_05226_),
    .C1(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__a211o_1 _12380_ (.A1(_05226_),
    .A2(_05227_),
    .B1(_05146_),
    .C1(_05147_),
    .X(_05229_));
 sky130_fd_sc_hd__o211ai_4 _12381_ (.A1(_05114_),
    .A2(_05145_),
    .B1(_05228_),
    .C1(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__a211o_1 _12382_ (.A1(_05228_),
    .A2(_05229_),
    .B1(_05114_),
    .C1(_05145_),
    .X(_05231_));
 sky130_fd_sc_hd__o211ai_4 _12383_ (.A1(_05120_),
    .A2(_05122_),
    .B1(_05230_),
    .C1(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__a211o_1 _12384_ (.A1(_05230_),
    .A2(_05231_),
    .B1(_05120_),
    .C1(_05122_),
    .X(_05233_));
 sky130_fd_sc_hd__or2_1 _12385_ (.A(_05087_),
    .B(_05089_),
    .X(_05234_));
 sky130_fd_sc_hd__o21ai_1 _12386_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__and3_1 _12387_ (.A(_05232_),
    .B(_05233_),
    .C(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__a21oi_1 _12388_ (.A1(_05232_),
    .A2(_05233_),
    .B1(_05235_),
    .Y(_05237_));
 sky130_fd_sc_hd__o211a_1 _12389_ (.A1(_05236_),
    .A2(_05237_),
    .B1(_05126_),
    .C1(_05128_),
    .X(_05238_));
 sky130_fd_sc_hd__a211oi_1 _12390_ (.A1(_05126_),
    .A2(_05128_),
    .B1(_05236_),
    .C1(_05237_),
    .Y(_05239_));
 sky130_fd_sc_hd__or2_1 _12391_ (.A(_05238_),
    .B(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__nor2_1 _12392_ (.A(_05130_),
    .B(_05131_),
    .Y(_05242_));
 sky130_fd_sc_hd__nor2_1 _12393_ (.A(_05242_),
    .B(_05136_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(_05240_),
    .B(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__o21a_1 _12395_ (.A1(_05240_),
    .A2(_05243_),
    .B1(_03133_),
    .X(_05245_));
 sky130_fd_sc_hd__xor2_1 _12396_ (.A(_02324_),
    .B(_02346_),
    .X(_05246_));
 sky130_fd_sc_hd__nor2_1 _12397_ (.A(_02398_),
    .B(_02584_),
    .Y(_05247_));
 sky130_fd_sc_hd__xnor2_2 _12398_ (.A(_05246_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__inv_2 _12399_ (.A(_02800_),
    .Y(_05249_));
 sky130_fd_sc_hd__a2bb2o_1 _12400_ (.A1_N(_04929_),
    .A2_N(_02727_),
    .B1(_05249_),
    .B2(_04011_),
    .X(_05250_));
 sky130_fd_sc_hd__a221o_1 _12401_ (.A1(\MuI.result[15] ),
    .A2(_02738_),
    .B1(_04642_),
    .B2(_04865_),
    .C1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__a32o_1 _12402_ (.A1(_02916_),
    .A2(_04929_),
    .A3(_02744_),
    .B1(_04627_),
    .B2(\FuI.Integer[15] ),
    .X(_05253_));
 sky130_fd_sc_hd__a221o_1 _12403_ (.A1(_04994_),
    .A2(_03675_),
    .B1(_02722_),
    .B2(_02916_),
    .C1(_05253_),
    .X(_05254_));
 sky130_fd_sc_hd__a21boi_1 _12404_ (.A1(_02795_),
    .A2(_05028_),
    .B1_N(_06629_),
    .Y(_05255_));
 sky130_fd_sc_hd__xnor2_1 _12405_ (.A(_05249_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__a22o_1 _12406_ (.A1(\AuI.result[15] ),
    .A2(_02938_),
    .B1(_05256_),
    .B2(_02935_),
    .X(_05257_));
 sky130_fd_sc_hd__or3_1 _12407_ (.A(_05251_),
    .B(_05254_),
    .C(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__a221o_1 _12408_ (.A1(_05244_),
    .A2(_05245_),
    .B1(_05248_),
    .B2(_03315_),
    .C1(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__a31o_4 _12409_ (.A1(_02752_),
    .A2(_05142_),
    .A3(_05143_),
    .B1(_05259_),
    .X(net75));
 sky130_fd_sc_hd__a21oi_1 _12410_ (.A1(_02796_),
    .A2(_02792_),
    .B1(_02799_),
    .Y(_05260_));
 sky130_fd_sc_hd__o31ai_1 _12411_ (.A1(_02795_),
    .A2(_05249_),
    .A3(_05017_),
    .B1(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(_05261_),
    .A1(_02899_),
    .S(_04635_),
    .X(_05263_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_02865_),
    .B(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(_02865_),
    .B(_05263_),
    .X(_05265_));
 sky130_fd_sc_hd__o211a_1 _12415_ (.A1(_05120_),
    .A2(_05122_),
    .B1(_05230_),
    .C1(_05231_),
    .X(_05266_));
 sky130_fd_sc_hd__and2_1 _12416_ (.A(_05149_),
    .B(_05157_),
    .X(_05267_));
 sky130_fd_sc_hd__or2_1 _12417_ (.A(_05041_),
    .B(_05151_),
    .X(_05268_));
 sky130_fd_sc_hd__xnor2_1 _12418_ (.A(_05154_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__a22oi_1 _12419_ (.A1(_01146_),
    .A2(_03425_),
    .B1(_03449_),
    .B2(_01147_),
    .Y(_05270_));
 sky130_fd_sc_hd__and4_1 _12420_ (.A(_00299_),
    .B(_00231_),
    .C(_00382_),
    .D(_06537_),
    .X(_05271_));
 sky130_fd_sc_hd__nor2_1 _12421_ (.A(_05270_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_1 _12422_ (.A(_00270_),
    .B(_03071_),
    .Y(_05274_));
 sky130_fd_sc_hd__xnor2_1 _12423_ (.A(_05272_),
    .B(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__a22oi_2 _12424_ (.A1(_03099_),
    .A2(_00785_),
    .B1(_05884_),
    .B2(_03056_),
    .Y(_05276_));
 sky130_fd_sc_hd__and4_1 _12425_ (.A(_00237_),
    .B(_00462_),
    .C(_00785_),
    .D(_00153_),
    .X(_05277_));
 sky130_fd_sc_hd__nand2_1 _12426_ (.A(_00088_),
    .B(_03247_),
    .Y(_05278_));
 sky130_fd_sc_hd__or3_1 _12427_ (.A(_05276_),
    .B(_05277_),
    .C(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__o21ai_1 _12428_ (.A1(_05276_),
    .A2(_05277_),
    .B1(_05278_),
    .Y(_05280_));
 sky130_fd_sc_hd__o21bai_1 _12429_ (.A1(_05164_),
    .A2(_05167_),
    .B1_N(_05165_),
    .Y(_05281_));
 sky130_fd_sc_hd__and3_1 _12430_ (.A(_05279_),
    .B(_05280_),
    .C(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__a21o_1 _12431_ (.A1(_05279_),
    .A2(_05280_),
    .B1(_05281_),
    .X(_05283_));
 sky130_fd_sc_hd__and2b_1 _12432_ (.A_N(_05282_),
    .B(_05283_),
    .X(_05285_));
 sky130_fd_sc_hd__xnor2_1 _12433_ (.A(_05275_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__or2_2 _12434_ (.A(_05269_),
    .B(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__nand2_1 _12435_ (.A(_05269_),
    .B(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__o211ai_4 _12436_ (.A1(_05267_),
    .A2(_05174_),
    .B1(_05287_),
    .C1(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__a211o_1 _12437_ (.A1(_05287_),
    .A2(_05288_),
    .B1(_05267_),
    .C1(_05174_),
    .X(_05290_));
 sky130_fd_sc_hd__or2b_1 _12438_ (.A(_05208_),
    .B_N(_05207_),
    .X(_05291_));
 sky130_fd_sc_hd__a22oi_1 _12439_ (.A1(_00676_),
    .A2(_06568_),
    .B1(_03047_),
    .B2(_00506_),
    .Y(_05292_));
 sky130_fd_sc_hd__and4_1 _12440_ (.A(_03539_),
    .B(_03593_),
    .C(_06518_),
    .D(_00412_),
    .X(_05293_));
 sky130_fd_sc_hd__nor2_1 _12441_ (.A(_05292_),
    .B(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand2_1 _12442_ (.A(_06439_),
    .B(_05198_),
    .Y(_05295_));
 sky130_fd_sc_hd__xnor2_1 _12443_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__o21ba_1 _12444_ (.A1(_05203_),
    .A2(_05206_),
    .B1_N(_05204_),
    .X(_05297_));
 sky130_fd_sc_hd__xnor2_1 _12445_ (.A(_05296_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand2_1 _12446_ (.A(_03722_),
    .B(_05123_),
    .Y(_05299_));
 sky130_fd_sc_hd__xor2_1 _12447_ (.A(_05298_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__a21o_1 _12448_ (.A1(_05291_),
    .A2(_05211_),
    .B1(_05300_),
    .X(_05301_));
 sky130_fd_sc_hd__nand3_1 _12449_ (.A(_05291_),
    .B(_05211_),
    .C(_05300_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_1 _12450_ (.A(_05301_),
    .B(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(net61),
    .B(_05058_),
    .Y(_05304_));
 sky130_fd_sc_hd__or2_1 _12452_ (.A(_05303_),
    .B(_05304_),
    .X(_05306_));
 sky130_fd_sc_hd__nand2_1 _12453_ (.A(_05303_),
    .B(_05304_),
    .Y(_05307_));
 sky130_fd_sc_hd__and2_1 _12454_ (.A(_05306_),
    .B(_05307_),
    .X(_05308_));
 sky130_fd_sc_hd__and2_1 _12455_ (.A(_05168_),
    .B(_05169_),
    .X(_05309_));
 sky130_fd_sc_hd__nand2_1 _12456_ (.A(_05188_),
    .B(_05190_),
    .Y(_05310_));
 sky130_fd_sc_hd__a31o_1 _12457_ (.A1(_00077_),
    .A2(_05520_),
    .A3(_05161_),
    .B1(_05160_),
    .X(_05311_));
 sky130_fd_sc_hd__a22oi_1 _12458_ (.A1(_00279_),
    .A2(_06666_),
    .B1(_00398_),
    .B2(_03378_),
    .Y(_05312_));
 sky130_fd_sc_hd__and4_1 _12459_ (.A(net113),
    .B(_03432_),
    .C(_06489_),
    .D(_05498_),
    .X(_05313_));
 sky130_fd_sc_hd__nor2_1 _12460_ (.A(_05312_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand2_1 _12461_ (.A(_00292_),
    .B(_06477_),
    .Y(_05315_));
 sky130_fd_sc_hd__xnor2_1 _12462_ (.A(_05314_),
    .B(_05315_),
    .Y(_05317_));
 sky130_fd_sc_hd__xor2_1 _12463_ (.A(_05311_),
    .B(_05317_),
    .X(_05318_));
 sky130_fd_sc_hd__xor2_1 _12464_ (.A(_05310_),
    .B(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__o21a_1 _12465_ (.A1(_05309_),
    .A2(_05171_),
    .B1(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__nor3_1 _12466_ (.A(_05309_),
    .B(_05171_),
    .C(_05319_),
    .Y(_05321_));
 sky130_fd_sc_hd__a211o_1 _12467_ (.A1(_05191_),
    .A2(_05195_),
    .B1(_05320_),
    .C1(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__o211ai_2 _12468_ (.A1(_05320_),
    .A2(_05321_),
    .B1(_05191_),
    .C1(_05195_),
    .Y(_05323_));
 sky130_fd_sc_hd__o211ai_1 _12469_ (.A1(_05196_),
    .A2(_05199_),
    .B1(_05322_),
    .C1(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__a211o_1 _12470_ (.A1(_05322_),
    .A2(_05323_),
    .B1(_05196_),
    .C1(_05199_),
    .X(_05325_));
 sky130_fd_sc_hd__and3_1 _12471_ (.A(_05308_),
    .B(_05324_),
    .C(_05325_),
    .X(_05326_));
 sky130_fd_sc_hd__a21oi_1 _12472_ (.A1(_05324_),
    .A2(_05325_),
    .B1(_05308_),
    .Y(_05328_));
 sky130_fd_sc_hd__or3_4 _12473_ (.A(_05178_),
    .B(_05326_),
    .C(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__o21ai_2 _12474_ (.A1(_05326_),
    .A2(_05328_),
    .B1(_05178_),
    .Y(_05330_));
 sky130_fd_sc_hd__o211ai_4 _12475_ (.A1(_05201_),
    .A2(_05219_),
    .B1(_05329_),
    .C1(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a211o_1 _12476_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05201_),
    .C1(_05219_),
    .X(_05332_));
 sky130_fd_sc_hd__and4_1 _12477_ (.A(_05289_),
    .B(_05290_),
    .C(_05331_),
    .D(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__a22oi_2 _12478_ (.A1(_05289_),
    .A2(_05290_),
    .B1(_05331_),
    .B2(_05332_),
    .Y(_05334_));
 sky130_fd_sc_hd__or3_4 _12479_ (.A(_05226_),
    .B(_05333_),
    .C(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__o21ai_2 _12480_ (.A1(_05333_),
    .A2(_05334_),
    .B1(_05226_),
    .Y(_05336_));
 sky130_fd_sc_hd__o211a_1 _12481_ (.A1(_05222_),
    .A2(_05224_),
    .B1(_05335_),
    .C1(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__a211oi_2 _12482_ (.A1(_05335_),
    .A2(_05336_),
    .B1(_05222_),
    .C1(_05224_),
    .Y(_05339_));
 sky130_fd_sc_hd__a211o_2 _12483_ (.A1(_05228_),
    .A2(_05230_),
    .B1(_05337_),
    .C1(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__o211ai_4 _12484_ (.A1(_05337_),
    .A2(_05339_),
    .B1(_05228_),
    .C1(_05230_),
    .Y(_05341_));
 sky130_fd_sc_hd__and2b_1 _12485_ (.A_N(_05213_),
    .B(_05215_),
    .X(_05342_));
 sky130_fd_sc_hd__a31o_1 _12486_ (.A1(_03842_),
    .A2(_04994_),
    .A3(_05216_),
    .B1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__nand3_1 _12487_ (.A(_05340_),
    .B(_05341_),
    .C(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__a21o_1 _12488_ (.A1(_05340_),
    .A2(_05341_),
    .B1(_05343_),
    .X(_05345_));
 sky130_fd_sc_hd__o211a_1 _12489_ (.A1(_05266_),
    .A2(_05236_),
    .B1(_05344_),
    .C1(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__a211oi_1 _12490_ (.A1(_05344_),
    .A2(_05345_),
    .B1(_05266_),
    .C1(_05236_),
    .Y(_05347_));
 sky130_fd_sc_hd__nor2_1 _12491_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__xor2_1 _12492_ (.A(_05130_),
    .B(_05131_),
    .X(_05350_));
 sky130_fd_sc_hd__nor2_1 _12493_ (.A(_05238_),
    .B(_05239_),
    .Y(_05351_));
 sky130_fd_sc_hd__and4bb_1 _12494_ (.A_N(_04872_),
    .B_N(_04998_),
    .C(_05350_),
    .D(_05351_),
    .X(_05352_));
 sky130_fd_sc_hd__inv_2 _12495_ (.A(_04997_),
    .Y(_05353_));
 sky130_fd_sc_hd__o2111a_1 _12496_ (.A1(_04999_),
    .A2(_04996_),
    .B1(_05353_),
    .C1(_05350_),
    .D1(_05351_),
    .X(_05354_));
 sky130_fd_sc_hd__o21ba_1 _12497_ (.A1(_05242_),
    .A2(_05239_),
    .B1_N(_05238_),
    .X(_05355_));
 sky130_fd_sc_hd__a211o_1 _12498_ (.A1(_04877_),
    .A2(_05352_),
    .B1(_05354_),
    .C1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__a21oi_1 _12499_ (.A1(_04873_),
    .A2(_05352_),
    .B1(_05356_),
    .Y(_05357_));
 sky130_fd_sc_hd__a211oi_2 _12500_ (.A1(_02703_),
    .A2(_04315_),
    .B1(_05356_),
    .C1(_04321_),
    .Y(_05358_));
 sky130_fd_sc_hd__nor2_1 _12501_ (.A(_05357_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__or2_1 _12502_ (.A(_05348_),
    .B(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__nand2_1 _12503_ (.A(_05348_),
    .B(_05359_),
    .Y(_05361_));
 sky130_fd_sc_hd__a2bb2o_1 _12504_ (.A1_N(_04994_),
    .A2_N(_02728_),
    .B1(_02732_),
    .B2(\AuI.result[16] ),
    .X(_05362_));
 sky130_fd_sc_hd__inv_2 _12505_ (.A(_02865_),
    .Y(_05363_));
 sky130_fd_sc_hd__a32o_1 _12506_ (.A1(_02970_),
    .A2(_04994_),
    .A3(_02743_),
    .B1(_02944_),
    .B2(_04929_),
    .X(_05364_));
 sky130_fd_sc_hd__a221o_1 _12507_ (.A1(\MuI.result[16] ),
    .A2(_02738_),
    .B1(_04011_),
    .B2(_05363_),
    .C1(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__a221o_1 _12508_ (.A1(\FuI.Integer[16] ),
    .A2(_02931_),
    .B1(_02719_),
    .B2(_05058_),
    .C1(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__a211o_1 _12509_ (.A1(_02970_),
    .A2(_02724_),
    .B1(_05362_),
    .C1(_05366_),
    .X(_05367_));
 sky130_fd_sc_hd__or2_1 _12510_ (.A(_02400_),
    .B(_02584_),
    .X(_05368_));
 sky130_fd_sc_hd__a21oi_2 _12511_ (.A1(_02621_),
    .A2(_05368_),
    .B1(_02619_),
    .Y(_05369_));
 sky130_fd_sc_hd__and3_1 _12512_ (.A(_02621_),
    .B(_05368_),
    .C(_02619_),
    .X(_05371_));
 sky130_fd_sc_hd__nand2_1 _12513_ (.A(_02916_),
    .B(_04929_),
    .Y(_05372_));
 sky130_fd_sc_hd__o21ai_1 _12514_ (.A1(_02800_),
    .A2(_05255_),
    .B1(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__nor2_1 _12515_ (.A(_05363_),
    .B(_05373_),
    .Y(_05374_));
 sky130_fd_sc_hd__and2_1 _12516_ (.A(_05363_),
    .B(_05373_),
    .X(_05375_));
 sky130_fd_sc_hd__or3_2 _12517_ (.A(_02711_),
    .B(_05374_),
    .C(_05375_),
    .X(_05376_));
 sky130_fd_sc_hd__o31ai_4 _12518_ (.A1(_04159_),
    .A2(_05369_),
    .A3(_05371_),
    .B1(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__a311o_1 _12519_ (.A1(_03134_),
    .A2(_05360_),
    .A3(_05361_),
    .B1(_05367_),
    .C1(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__a31o_4 _12520_ (.A1(_02752_),
    .A2(_05264_),
    .A3(_05265_),
    .B1(_05378_),
    .X(net76));
 sky130_fd_sc_hd__inv_2 _12521_ (.A(_02849_),
    .Y(_05379_));
 sky130_fd_sc_hd__nor2_1 _12522_ (.A(_05379_),
    .B(_02850_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21o_1 _12523_ (.A1(_02865_),
    .A2(_05261_),
    .B1(_02864_),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _12524_ (.A0(_05382_),
    .A1(_02900_),
    .S(_04635_),
    .X(_05383_));
 sky130_fd_sc_hd__nand2_1 _12525_ (.A(_05381_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__or2_1 _12526_ (.A(_05381_),
    .B(_05383_),
    .X(_05385_));
 sky130_fd_sc_hd__a32o_1 _12527_ (.A1(_02621_),
    .A2(_05368_),
    .A3(_02619_),
    .B1(_02618_),
    .B2(_02617_),
    .X(_05386_));
 sky130_fd_sc_hd__xor2_2 _12528_ (.A(_02613_),
    .B(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a21oi_1 _12529_ (.A1(_02970_),
    .A2(_04994_),
    .B1(_05375_),
    .Y(_05388_));
 sky130_fd_sc_hd__xnor2_1 _12530_ (.A(_02853_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a22o_1 _12531_ (.A1(_03024_),
    .A2(_02721_),
    .B1(_02853_),
    .B2(_04011_),
    .X(_05390_));
 sky130_fd_sc_hd__a221o_1 _12532_ (.A1(\MuI.result[17] ),
    .A2(_02738_),
    .B1(_02931_),
    .B2(\FuI.Integer[17] ),
    .C1(_05390_),
    .X(_05392_));
 sky130_fd_sc_hd__nor2_1 _12533_ (.A(_05058_),
    .B(_02727_),
    .Y(_05393_));
 sky130_fd_sc_hd__a31o_1 _12534_ (.A1(_03024_),
    .A2(_05058_),
    .A3(_02744_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__a221o_1 _12535_ (.A1(_05134_),
    .A2(_03675_),
    .B1(_04642_),
    .B2(_04994_),
    .C1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__a211o_1 _12536_ (.A1(\AuI.result[17] ),
    .A2(_02732_),
    .B1(_05392_),
    .C1(_05395_),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _12537_ (.A1(_03489_),
    .A2(_05389_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__o211ai_4 _12538_ (.A1(_05222_),
    .A2(_05224_),
    .B1(_05335_),
    .C1(_05336_),
    .Y(_05398_));
 sky130_fd_sc_hd__or2_1 _12539_ (.A(_05154_),
    .B(_05268_),
    .X(_05399_));
 sky130_fd_sc_hd__a22oi_1 _12540_ (.A1(_03282_),
    .A2(_05702_),
    .B1(_05767_),
    .B2(_03228_),
    .Y(_05400_));
 sky130_fd_sc_hd__and4_1 _12541_ (.A(_00299_),
    .B(_00231_),
    .C(_06537_),
    .D(_00385_),
    .X(_05401_));
 sky130_fd_sc_hd__nor2_1 _12542_ (.A(_05400_),
    .B(_05401_),
    .Y(_05403_));
 sky130_fd_sc_hd__nand2_1 _12543_ (.A(_00270_),
    .B(_05649_),
    .Y(_05404_));
 sky130_fd_sc_hd__xnor2_1 _12544_ (.A(_05403_),
    .B(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__a22o_1 _12545_ (.A1(_00081_),
    .A2(_03082_),
    .B1(_00789_),
    .B2(_00086_),
    .X(_05406_));
 sky130_fd_sc_hd__nand4_1 _12546_ (.A(_00133_),
    .B(_00132_),
    .C(_05884_),
    .D(_00789_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand4_1 _12547_ (.A(_03174_),
    .B(_03257_),
    .C(_05406_),
    .D(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__a22o_1 _12548_ (.A1(_00262_),
    .A2(_03257_),
    .B1(_05406_),
    .B2(_05407_),
    .X(_05409_));
 sky130_fd_sc_hd__o21bai_1 _12549_ (.A1(_05276_),
    .A2(_05278_),
    .B1_N(_05277_),
    .Y(_05410_));
 sky130_fd_sc_hd__and3_1 _12550_ (.A(_05408_),
    .B(_05409_),
    .C(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__a21o_1 _12551_ (.A1(_05408_),
    .A2(_05409_),
    .B1(_05410_),
    .X(_05412_));
 sky130_fd_sc_hd__or2b_1 _12552_ (.A(_05411_),
    .B_N(_05412_),
    .X(_05414_));
 sky130_fd_sc_hd__xor2_1 _12553_ (.A(_05405_),
    .B(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__or3_1 _12554_ (.A(_05039_),
    .B(_05151_),
    .C(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__o21ai_1 _12555_ (.A1(_05039_),
    .A2(_05151_),
    .B1(_05415_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _12556_ (.A(_05416_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21o_1 _12557_ (.A1(_05399_),
    .A2(_05287_),
    .B1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__nand3_1 _12558_ (.A(_05399_),
    .B(_05287_),
    .C(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_1 _12559_ (.A(_05419_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__o211a_1 _12560_ (.A1(_05196_),
    .A2(_05199_),
    .B1(_05322_),
    .C1(_05323_),
    .X(_05422_));
 sky130_fd_sc_hd__or2b_1 _12561_ (.A(_05297_),
    .B_N(_05296_),
    .X(_05423_));
 sky130_fd_sc_hd__nand3_1 _12562_ (.A(_03733_),
    .B(_05123_),
    .C(_05298_),
    .Y(_05424_));
 sky130_fd_sc_hd__a22oi_1 _12563_ (.A1(_00676_),
    .A2(_03047_),
    .B1(_06477_),
    .B2(_06444_),
    .Y(_05425_));
 sky130_fd_sc_hd__and4_1 _12564_ (.A(_06434_),
    .B(_00678_),
    .C(_00412_),
    .D(_00530_),
    .X(_05426_));
 sky130_fd_sc_hd__nor2_1 _12565_ (.A(_05425_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_03658_),
    .B(_05262_),
    .Y(_05428_));
 sky130_fd_sc_hd__xnor2_1 _12567_ (.A(_05427_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__a31o_1 _12568_ (.A1(_03525_),
    .A2(_05198_),
    .A3(_05294_),
    .B1(_05293_),
    .X(_05430_));
 sky130_fd_sc_hd__xor2_1 _12569_ (.A(_05429_),
    .B(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__and2_1 _12570_ (.A(_03722_),
    .B(_05209_),
    .X(_05432_));
 sky130_fd_sc_hd__xnor2_1 _12571_ (.A(_05431_),
    .B(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__a21oi_2 _12572_ (.A1(_05423_),
    .A2(_05424_),
    .B1(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__and3_1 _12573_ (.A(_05423_),
    .B(_05424_),
    .C(_05433_),
    .X(_05436_));
 sky130_fd_sc_hd__nor2_1 _12574_ (.A(_05435_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__nand2_1 _12575_ (.A(_00502_),
    .B(_05123_),
    .Y(_05438_));
 sky130_fd_sc_hd__xnor2_1 _12576_ (.A(_05437_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_1 _12577_ (.A1(_05309_),
    .A2(_05171_),
    .B1(_05319_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _12578_ (.A(_05311_),
    .B(_05317_),
    .Y(_05441_));
 sky130_fd_sc_hd__nand2_1 _12579_ (.A(_05310_),
    .B(_05318_),
    .Y(_05442_));
 sky130_fd_sc_hd__a21o_1 _12580_ (.A1(_05275_),
    .A2(_05283_),
    .B1(_05282_),
    .X(_05443_));
 sky130_fd_sc_hd__a31o_1 _12581_ (.A1(_03497_),
    .A2(_05391_),
    .A3(_05314_),
    .B1(_05313_),
    .X(_05444_));
 sky130_fd_sc_hd__o21bai_1 _12582_ (.A1(_05270_),
    .A2(_05274_),
    .B1_N(_05271_),
    .Y(_05446_));
 sky130_fd_sc_hd__a22o_1 _12583_ (.A1(_00289_),
    .A2(_00398_),
    .B1(_03424_),
    .B2(_03378_),
    .X(_05447_));
 sky130_fd_sc_hd__nand4_2 _12584_ (.A(_00290_),
    .B(_00289_),
    .C(_05509_),
    .D(_03424_),
    .Y(_05448_));
 sky130_fd_sc_hd__a22o_1 _12585_ (.A1(_00283_),
    .A2(_06546_),
    .B1(_05447_),
    .B2(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__nand4_2 _12586_ (.A(_03486_),
    .B(_05456_),
    .C(_05447_),
    .D(_05448_),
    .Y(_05450_));
 sky130_fd_sc_hd__nand3_2 _12587_ (.A(_05446_),
    .B(_05449_),
    .C(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__a21o_1 _12588_ (.A1(_05449_),
    .A2(_05450_),
    .B1(_05446_),
    .X(_05452_));
 sky130_fd_sc_hd__nand3_2 _12589_ (.A(_05444_),
    .B(_05451_),
    .C(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__a21o_1 _12590_ (.A1(_05451_),
    .A2(_05452_),
    .B1(_05444_),
    .X(_05454_));
 sky130_fd_sc_hd__and3_2 _12591_ (.A(_05443_),
    .B(_05453_),
    .C(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__a21oi_2 _12592_ (.A1(_05453_),
    .A2(_05454_),
    .B1(_05443_),
    .Y(_05457_));
 sky130_fd_sc_hd__a211oi_4 _12593_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05455_),
    .C1(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__o211a_1 _12594_ (.A1(_05455_),
    .A2(_05457_),
    .B1(_05441_),
    .C1(_05442_),
    .X(_05459_));
 sky130_fd_sc_hd__a211o_1 _12595_ (.A1(_05440_),
    .A2(_05322_),
    .B1(_05458_),
    .C1(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__o211ai_1 _12596_ (.A1(_05458_),
    .A2(_05459_),
    .B1(_05440_),
    .C1(_05322_),
    .Y(_05461_));
 sky130_fd_sc_hd__and3_1 _12597_ (.A(_05439_),
    .B(_05460_),
    .C(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__a21oi_1 _12598_ (.A1(_05460_),
    .A2(_05461_),
    .B1(_05439_),
    .Y(_05463_));
 sky130_fd_sc_hd__or3_1 _12599_ (.A(_05289_),
    .B(_05462_),
    .C(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__o21ai_1 _12600_ (.A1(_05462_),
    .A2(_05463_),
    .B1(_05289_),
    .Y(_05465_));
 sky130_fd_sc_hd__o211a_1 _12601_ (.A1(_05422_),
    .A2(_05326_),
    .B1(_05464_),
    .C1(_05465_),
    .X(_05466_));
 sky130_fd_sc_hd__a211oi_1 _12602_ (.A1(_05464_),
    .A2(_05465_),
    .B1(_05422_),
    .C1(_05326_),
    .Y(_05468_));
 sky130_fd_sc_hd__or3_2 _12603_ (.A(_05421_),
    .B(_05466_),
    .C(_05468_),
    .X(_05469_));
 sky130_fd_sc_hd__o21ai_1 _12604_ (.A1(_05466_),
    .A2(_05468_),
    .B1(_05421_),
    .Y(_05470_));
 sky130_fd_sc_hd__and3_2 _12605_ (.A(_05333_),
    .B(_05469_),
    .C(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__a21oi_2 _12606_ (.A1(_05469_),
    .A2(_05470_),
    .B1(_05333_),
    .Y(_05472_));
 sky130_fd_sc_hd__a211oi_4 _12607_ (.A1(_05329_),
    .A2(_05331_),
    .B1(_05471_),
    .C1(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__o211a_1 _12608_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05329_),
    .C1(_05331_),
    .X(_05474_));
 sky130_fd_sc_hd__a211oi_4 _12609_ (.A1(_05335_),
    .A2(_05398_),
    .B1(_05473_),
    .C1(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__o211a_1 _12610_ (.A1(_05473_),
    .A2(_05474_),
    .B1(_05335_),
    .C1(_05398_),
    .X(_05476_));
 sky130_fd_sc_hd__a211oi_2 _12611_ (.A1(_05301_),
    .A2(_05306_),
    .B1(_05475_),
    .C1(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__o211a_1 _12612_ (.A1(_05475_),
    .A2(_05476_),
    .B1(_05301_),
    .C1(_05306_),
    .X(_05479_));
 sky130_fd_sc_hd__a211oi_1 _12613_ (.A1(_05340_),
    .A2(_05344_),
    .B1(_05477_),
    .C1(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__o211ai_1 _12614_ (.A1(_05477_),
    .A2(_05479_),
    .B1(_05340_),
    .C1(_05344_),
    .Y(_05481_));
 sky130_fd_sc_hd__and2b_1 _12615_ (.A_N(_05480_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__a21o_1 _12616_ (.A1(_05348_),
    .A2(_05359_),
    .B1(_05346_),
    .X(_05483_));
 sky130_fd_sc_hd__a21oi_1 _12617_ (.A1(_05482_),
    .A2(_05483_),
    .B1(_06427_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21a_1 _12618_ (.A1(_05482_),
    .A2(_05483_),
    .B1(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__a211o_1 _12619_ (.A1(_03315_),
    .A2(_05387_),
    .B1(_05397_),
    .C1(_05485_),
    .X(_05486_));
 sky130_fd_sc_hd__a31o_2 _12620_ (.A1(_02752_),
    .A2(_05384_),
    .A3(_05385_),
    .B1(_05486_),
    .X(net77));
 sky130_fd_sc_hd__a21o_1 _12621_ (.A1(_02852_),
    .A2(_05382_),
    .B1(_05379_),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_1 _12622_ (.A0(_05487_),
    .A1(_02901_),
    .S(_02928_),
    .X(_05488_));
 sky130_fd_sc_hd__or2_1 _12623_ (.A(_02856_),
    .B(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__nand2_1 _12624_ (.A(_02856_),
    .B(_05488_),
    .Y(_05490_));
 sky130_fd_sc_hd__and3_1 _12625_ (.A(_03831_),
    .B(_05134_),
    .C(_05437_),
    .X(_05491_));
 sky130_fd_sc_hd__nor3_2 _12626_ (.A(_05289_),
    .B(_05462_),
    .C(_05463_),
    .Y(_05492_));
 sky130_fd_sc_hd__and4_1 _12627_ (.A(_00921_),
    .B(_01206_),
    .C(_03444_),
    .D(_05948_),
    .X(_05493_));
 sky130_fd_sc_hd__and4_1 _12628_ (.A(_00262_),
    .B(_03257_),
    .C(_05406_),
    .D(_05407_),
    .X(_05494_));
 sky130_fd_sc_hd__a22o_1 _12629_ (.A1(_00262_),
    .A2(_05895_),
    .B1(_05959_),
    .B2(_03110_),
    .X(_05495_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(_01206_),
    .B(_03444_),
    .Y(_05496_));
 sky130_fd_sc_hd__or3_1 _12631_ (.A(_02801_),
    .B(_02875_),
    .C(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__o211a_1 _12632_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_05495_),
    .C1(_05497_),
    .X(_05499_));
 sky130_fd_sc_hd__a211o_1 _12633_ (.A1(_05495_),
    .A2(_05497_),
    .B1(_05493_),
    .C1(_05494_),
    .X(_05500_));
 sky130_fd_sc_hd__and2b_1 _12634_ (.A_N(_05499_),
    .B(_05500_),
    .X(_05501_));
 sky130_fd_sc_hd__a22oi_1 _12635_ (.A1(_01146_),
    .A2(_03247_),
    .B1(_05820_),
    .B2(_03228_),
    .Y(_05502_));
 sky130_fd_sc_hd__and4_1 _12636_ (.A(_00299_),
    .B(_00231_),
    .C(_00385_),
    .D(_00783_),
    .X(_05503_));
 sky130_fd_sc_hd__nor2_1 _12637_ (.A(_05502_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2_1 _12638_ (.A(_00270_),
    .B(_03449_),
    .Y(_05505_));
 sky130_fd_sc_hd__xnor2_1 _12639_ (.A(_05504_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__xnor2_1 _12640_ (.A(_05501_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__or2_1 _12641_ (.A(_05416_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__nand2_1 _12642_ (.A(_05416_),
    .B(_05507_),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _12643_ (.A(_05508_),
    .B(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__a211oi_1 _12644_ (.A1(_05440_),
    .A2(_05322_),
    .B1(_05458_),
    .C1(_05459_),
    .Y(_05512_));
 sky130_fd_sc_hd__a22oi_1 _12645_ (.A1(_00676_),
    .A2(_05380_),
    .B1(_05445_),
    .B2(_00506_),
    .Y(_05513_));
 sky130_fd_sc_hd__and4_1 _12646_ (.A(_06434_),
    .B(_00678_),
    .C(_00530_),
    .D(_06666_),
    .X(_05514_));
 sky130_fd_sc_hd__nor2_1 _12647_ (.A(_05513_),
    .B(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__nand2_1 _12648_ (.A(_06439_),
    .B(_05327_),
    .Y(_05516_));
 sky130_fd_sc_hd__xnor2_1 _12649_ (.A(_05515_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__a31o_1 _12650_ (.A1(_02965_),
    .A2(_05262_),
    .A3(_05427_),
    .B1(_05426_),
    .X(_05518_));
 sky130_fd_sc_hd__xor2_1 _12651_ (.A(_05517_),
    .B(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__and2_1 _12652_ (.A(net60),
    .B(_05262_),
    .X(_05521_));
 sky130_fd_sc_hd__xnor2_1 _12653_ (.A(_05519_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__and2_1 _12654_ (.A(_05429_),
    .B(_05430_),
    .X(_05523_));
 sky130_fd_sc_hd__a21oi_1 _12655_ (.A1(_05431_),
    .A2(_05432_),
    .B1(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__xnor2_1 _12656_ (.A(_05522_),
    .B(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _12657_ (.A(net61),
    .B(_05209_),
    .Y(_05526_));
 sky130_fd_sc_hd__xor2_1 _12658_ (.A(_05525_),
    .B(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__a21o_1 _12659_ (.A1(_05405_),
    .A2(_05412_),
    .B1(_05411_),
    .X(_05528_));
 sky130_fd_sc_hd__o21bai_1 _12660_ (.A1(_05400_),
    .A2(_05404_),
    .B1_N(_05401_),
    .Y(_05529_));
 sky130_fd_sc_hd__a22o_1 _12661_ (.A1(_00279_),
    .A2(_03424_),
    .B1(_00382_),
    .B2(_00278_),
    .X(_05530_));
 sky130_fd_sc_hd__nand4_1 _12662_ (.A(_03378_),
    .B(_00289_),
    .C(_03424_),
    .D(_00382_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand4_1 _12663_ (.A(_03486_),
    .B(_05520_),
    .C(_05530_),
    .D(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__a22o_1 _12664_ (.A1(_00292_),
    .A2(_03051_),
    .B1(_05530_),
    .B2(_05532_),
    .X(_05534_));
 sky130_fd_sc_hd__nand3_1 _12665_ (.A(_05529_),
    .B(_05533_),
    .C(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__a21o_1 _12666_ (.A1(_05533_),
    .A2(_05534_),
    .B1(_05529_),
    .X(_05536_));
 sky130_fd_sc_hd__nand2_1 _12667_ (.A(_05448_),
    .B(_05450_),
    .Y(_05537_));
 sky130_fd_sc_hd__a21o_1 _12668_ (.A1(_05535_),
    .A2(_05536_),
    .B1(_05537_),
    .X(_05538_));
 sky130_fd_sc_hd__nand3_1 _12669_ (.A(_05537_),
    .B(_05535_),
    .C(_05536_),
    .Y(_05539_));
 sky130_fd_sc_hd__and3_1 _12670_ (.A(_05528_),
    .B(_05538_),
    .C(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__a21oi_1 _12671_ (.A1(_05538_),
    .A2(_05539_),
    .B1(_05528_),
    .Y(_05541_));
 sky130_fd_sc_hd__a211o_1 _12672_ (.A1(_05451_),
    .A2(_05453_),
    .B1(_05540_),
    .C1(_05541_),
    .X(_05543_));
 sky130_fd_sc_hd__o211ai_1 _12673_ (.A1(_05540_),
    .A2(_05541_),
    .B1(_05451_),
    .C1(_05453_),
    .Y(_05544_));
 sky130_fd_sc_hd__o211ai_2 _12674_ (.A1(_05455_),
    .A2(_05458_),
    .B1(_05543_),
    .C1(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__a211o_1 _12675_ (.A1(_05543_),
    .A2(_05544_),
    .B1(_05455_),
    .C1(_05458_),
    .X(_05546_));
 sky130_fd_sc_hd__and3_1 _12676_ (.A(_05527_),
    .B(_05545_),
    .C(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__a21oi_1 _12677_ (.A1(_05545_),
    .A2(_05546_),
    .B1(_05527_),
    .Y(_05548_));
 sky130_fd_sc_hd__or3_1 _12678_ (.A(_05419_),
    .B(_05547_),
    .C(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__o21ai_1 _12679_ (.A1(_05547_),
    .A2(_05548_),
    .B1(_05419_),
    .Y(_05550_));
 sky130_fd_sc_hd__o211a_1 _12680_ (.A1(_05512_),
    .A2(_05462_),
    .B1(_05549_),
    .C1(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__a211oi_1 _12681_ (.A1(_05549_),
    .A2(_05550_),
    .B1(_05512_),
    .C1(_05462_),
    .Y(_05552_));
 sky130_fd_sc_hd__nor3_2 _12682_ (.A(_05511_),
    .B(_05551_),
    .C(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21a_1 _12683_ (.A1(_05551_),
    .A2(_05552_),
    .B1(_05511_),
    .X(_05554_));
 sky130_fd_sc_hd__or3_4 _12684_ (.A(_05469_),
    .B(_05553_),
    .C(_05554_),
    .X(_05555_));
 sky130_fd_sc_hd__o21ai_2 _12685_ (.A1(_05553_),
    .A2(_05554_),
    .B1(_05469_),
    .Y(_05556_));
 sky130_fd_sc_hd__o211ai_4 _12686_ (.A1(_05492_),
    .A2(_05466_),
    .B1(_05555_),
    .C1(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__a211o_1 _12687_ (.A1(_05555_),
    .A2(_05556_),
    .B1(_05492_),
    .C1(_05466_),
    .X(_05558_));
 sky130_fd_sc_hd__o211ai_4 _12688_ (.A1(_05471_),
    .A2(_05473_),
    .B1(_05557_),
    .C1(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__a211o_1 _12689_ (.A1(_05557_),
    .A2(_05558_),
    .B1(_05471_),
    .C1(_05473_),
    .X(_05560_));
 sky130_fd_sc_hd__o211ai_2 _12690_ (.A1(_05435_),
    .A2(_05491_),
    .B1(_05559_),
    .C1(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__a211o_1 _12691_ (.A1(_05559_),
    .A2(_05560_),
    .B1(_05435_),
    .C1(_05491_),
    .X(_05562_));
 sky130_fd_sc_hd__and2_1 _12692_ (.A(_05561_),
    .B(_05562_),
    .X(_05564_));
 sky130_fd_sc_hd__o21ai_1 _12693_ (.A1(_05475_),
    .A2(_05477_),
    .B1(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__or3_1 _12694_ (.A(_05475_),
    .B(_05477_),
    .C(_05564_),
    .X(_05566_));
 sky130_fd_sc_hd__and2_1 _12695_ (.A(_05565_),
    .B(_05566_),
    .X(_05567_));
 sky130_fd_sc_hd__o21a_1 _12696_ (.A1(_05346_),
    .A2(_05480_),
    .B1(_05481_),
    .X(_05568_));
 sky130_fd_sc_hd__a31o_1 _12697_ (.A1(_05348_),
    .A2(_05359_),
    .A3(_05482_),
    .B1(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__nand2_1 _12698_ (.A(_05567_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21a_1 _12699_ (.A1(_05567_),
    .A2(_05569_),
    .B1(_03133_),
    .X(_05571_));
 sky130_fd_sc_hd__nand2_1 _12700_ (.A(_02613_),
    .B(_05386_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_02607_),
    .B(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(_02614_),
    .B(_02609_),
    .X(_05575_));
 sky130_fd_sc_hd__a21o_1 _12703_ (.A1(_05575_),
    .A2(_05572_),
    .B1(_02607_),
    .X(_05576_));
 sky130_fd_sc_hd__o211a_2 _12704_ (.A1(_02623_),
    .A2(_05573_),
    .B1(_05576_),
    .C1(_03314_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_1 _12705_ (.A(_02970_),
    .B(_04994_),
    .Y(_05578_));
 sky130_fd_sc_hd__nor2_1 _12706_ (.A(_03024_),
    .B(_05058_),
    .Y(_05579_));
 sky130_fd_sc_hd__a21oi_1 _12707_ (.A1(_05578_),
    .A2(_03186_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a31o_1 _12708_ (.A1(_05363_),
    .A2(_02853_),
    .A3(_05373_),
    .B1(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__or2b_1 _12709_ (.A(_02856_),
    .B_N(_05581_),
    .X(_05582_));
 sky130_fd_sc_hd__or2b_1 _12710_ (.A(_05581_),
    .B_N(_02856_),
    .X(_05583_));
 sky130_fd_sc_hd__o211ai_1 _12711_ (.A1(_02129_),
    .A2(_02854_),
    .B1(_02855_),
    .C1(_04011_),
    .Y(_05584_));
 sky130_fd_sc_hd__o21ai_1 _12712_ (.A1(_05134_),
    .A2(_02728_),
    .B1(_05584_),
    .Y(_05586_));
 sky130_fd_sc_hd__a22o_1 _12713_ (.A1(_02744_),
    .A2(_03974_),
    .B1(_02944_),
    .B2(_05058_),
    .X(_05587_));
 sky130_fd_sc_hd__a22o_1 _12714_ (.A1(\FuI.Integer[18] ),
    .A2(_06045_),
    .B1(_02718_),
    .B2(_05209_),
    .X(_05588_));
 sky130_fd_sc_hd__a211o_1 _12715_ (.A1(\MuI.result[18] ),
    .A2(_02738_),
    .B1(_05587_),
    .C1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__a211o_1 _12716_ (.A1(\AuI.result[18] ),
    .A2(_02732_),
    .B1(_05586_),
    .C1(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__a31o_1 _12717_ (.A1(_03489_),
    .A2(_05582_),
    .A3(_05583_),
    .B1(_05590_),
    .X(_05591_));
 sky130_fd_sc_hd__a211o_1 _12718_ (.A1(_05570_),
    .A2(_05571_),
    .B1(_05577_),
    .C1(_05591_),
    .X(_05592_));
 sky130_fd_sc_hd__a31o_4 _12719_ (.A1(_02752_),
    .A2(_05489_),
    .A3(_05490_),
    .B1(_05592_),
    .X(net78));
 sky130_fd_sc_hd__and2b_1 _12720_ (.A_N(_05134_),
    .B(_03067_),
    .X(_05593_));
 sky130_fd_sc_hd__a21o_1 _12721_ (.A1(_02856_),
    .A2(_05487_),
    .B1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_05594_),
    .A1(_02903_),
    .S(_02925_),
    .X(_05596_));
 sky130_fd_sc_hd__nand2_1 _12723_ (.A(_02868_),
    .B(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__o211a_1 _12724_ (.A1(_02868_),
    .A2(_05596_),
    .B1(_05597_),
    .C1(_02750_),
    .X(_05598_));
 sky130_fd_sc_hd__or2_1 _12725_ (.A(_05522_),
    .B(_05524_),
    .X(_05599_));
 sky130_fd_sc_hd__or2_1 _12726_ (.A(_05525_),
    .B(_05526_),
    .X(_05600_));
 sky130_fd_sc_hd__inv_2 _12727_ (.A(_05551_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_1 _12728_ (.A(_03228_),
    .B(_05820_),
    .Y(_05602_));
 sky130_fd_sc_hd__nand2_1 _12729_ (.A(_00125_),
    .B(_05884_),
    .Y(_05603_));
 sky130_fd_sc_hd__a22o_1 _12730_ (.A1(_00231_),
    .A2(_00785_),
    .B1(_05884_),
    .B2(_00299_),
    .X(_05604_));
 sky130_fd_sc_hd__o21ai_1 _12731_ (.A1(_05602_),
    .A2(_05603_),
    .B1(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__and2_1 _12732_ (.A(net114),
    .B(_00385_),
    .X(_05607_));
 sky130_fd_sc_hd__xnor2_1 _12733_ (.A(_05605_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__and3_1 _12734_ (.A(_03174_),
    .B(_05970_),
    .C(_05496_),
    .X(_05609_));
 sky130_fd_sc_hd__xnor2_1 _12735_ (.A(_05608_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__inv_2 _12736_ (.A(_05547_),
    .Y(_05611_));
 sky130_fd_sc_hd__a211oi_1 _12737_ (.A1(_05451_),
    .A2(_05453_),
    .B1(_05540_),
    .C1(_05541_),
    .Y(_05612_));
 sky130_fd_sc_hd__a21o_1 _12738_ (.A1(_05500_),
    .A2(_05506_),
    .B1(_05499_),
    .X(_05613_));
 sky130_fd_sc_hd__nand2_1 _12739_ (.A(_05532_),
    .B(_05533_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21bai_1 _12740_ (.A1(_05502_),
    .A2(_05505_),
    .B1_N(_05503_),
    .Y(_05615_));
 sky130_fd_sc_hd__a22o_1 _12741_ (.A1(_00279_),
    .A2(_00382_),
    .B1(_00163_),
    .B2(_03378_),
    .X(_05616_));
 sky130_fd_sc_hd__nand4_1 _12742_ (.A(_00290_),
    .B(_00289_),
    .C(_03425_),
    .D(_00163_),
    .Y(_05617_));
 sky130_fd_sc_hd__a22o_1 _12743_ (.A1(_00283_),
    .A2(_03071_),
    .B1(_05616_),
    .B2(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__nand4_1 _12744_ (.A(_03486_),
    .B(_05585_),
    .C(_05616_),
    .D(_05617_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand3_1 _12745_ (.A(_05615_),
    .B(_05618_),
    .C(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__a21o_1 _12746_ (.A1(_05618_),
    .A2(_05619_),
    .B1(_05615_),
    .X(_05621_));
 sky130_fd_sc_hd__nand3_1 _12747_ (.A(_05614_),
    .B(_05620_),
    .C(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__a21o_1 _12748_ (.A1(_05620_),
    .A2(_05621_),
    .B1(_05614_),
    .X(_05623_));
 sky130_fd_sc_hd__and3_1 _12749_ (.A(_05613_),
    .B(_05622_),
    .C(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__a21oi_1 _12750_ (.A1(_05622_),
    .A2(_05623_),
    .B1(_05613_),
    .Y(_05625_));
 sky130_fd_sc_hd__a211o_1 _12751_ (.A1(_05535_),
    .A2(_05539_),
    .B1(_05624_),
    .C1(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__o211ai_1 _12752_ (.A1(_05624_),
    .A2(_05625_),
    .B1(_05535_),
    .C1(_05539_),
    .Y(_05628_));
 sky130_fd_sc_hd__o211a_1 _12753_ (.A1(_05540_),
    .A2(_05612_),
    .B1(_05626_),
    .C1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__a211oi_1 _12754_ (.A1(_05626_),
    .A2(_05628_),
    .B1(_05540_),
    .C1(_05612_),
    .Y(_05630_));
 sky130_fd_sc_hd__a22oi_1 _12755_ (.A1(_00676_),
    .A2(_05445_),
    .B1(_05509_),
    .B2(_00506_),
    .Y(_05631_));
 sky130_fd_sc_hd__and4_1 _12756_ (.A(_03539_),
    .B(_00678_),
    .C(_06666_),
    .D(_00398_),
    .X(_05632_));
 sky130_fd_sc_hd__nor2_1 _12757_ (.A(_05631_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_1 _12758_ (.A(_06439_),
    .B(_05391_),
    .Y(_05634_));
 sky130_fd_sc_hd__xnor2_1 _12759_ (.A(_05633_),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ba_1 _12760_ (.A1(_05513_),
    .A2(_05516_),
    .B1_N(_05514_),
    .X(_05636_));
 sky130_fd_sc_hd__xnor2_1 _12761_ (.A(_05635_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _12762_ (.A(_06429_),
    .B(_05327_),
    .Y(_05639_));
 sky130_fd_sc_hd__xor2_1 _12763_ (.A(_05637_),
    .B(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__and2_1 _12764_ (.A(_05517_),
    .B(_05518_),
    .X(_05641_));
 sky130_fd_sc_hd__a21o_1 _12765_ (.A1(_05519_),
    .A2(_05521_),
    .B1(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__xnor2_1 _12766_ (.A(_05640_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2_1 _12767_ (.A(net61),
    .B(_05262_),
    .Y(_05644_));
 sky130_fd_sc_hd__xnor2_1 _12768_ (.A(_05643_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__nor3b_1 _12769_ (.A(_05629_),
    .B(_05630_),
    .C_N(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__o21ba_1 _12770_ (.A1(_05629_),
    .A2(_05630_),
    .B1_N(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__nor3_2 _12771_ (.A(_05508_),
    .B(_05646_),
    .C(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21a_1 _12772_ (.A1(_05646_),
    .A2(_05647_),
    .B1(_05508_),
    .X(_05650_));
 sky130_fd_sc_hd__a211oi_2 _12773_ (.A1(_05545_),
    .A2(_05611_),
    .B1(_05648_),
    .C1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__o211a_1 _12774_ (.A1(_05648_),
    .A2(_05650_),
    .B1(_05545_),
    .C1(_05611_),
    .X(_05652_));
 sky130_fd_sc_hd__or3_1 _12775_ (.A(_05610_),
    .B(_05651_),
    .C(_05652_),
    .X(_05653_));
 sky130_fd_sc_hd__o21ai_1 _12776_ (.A1(_05651_),
    .A2(_05652_),
    .B1(_05610_),
    .Y(_05654_));
 sky130_fd_sc_hd__and3_1 _12777_ (.A(_05553_),
    .B(_05653_),
    .C(_05654_),
    .X(_05655_));
 sky130_fd_sc_hd__a21oi_1 _12778_ (.A1(_05653_),
    .A2(_05654_),
    .B1(_05553_),
    .Y(_05656_));
 sky130_fd_sc_hd__or2_1 _12779_ (.A(_05655_),
    .B(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__a21oi_2 _12780_ (.A1(_05549_),
    .A2(_05601_),
    .B1(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__and3_1 _12781_ (.A(_05549_),
    .B(_05601_),
    .C(_05657_),
    .X(_05659_));
 sky130_fd_sc_hd__a211oi_4 _12782_ (.A1(_05555_),
    .A2(_05557_),
    .B1(_05658_),
    .C1(_05659_),
    .Y(_05661_));
 sky130_fd_sc_hd__o211a_1 _12783_ (.A1(_05658_),
    .A2(_05659_),
    .B1(_05555_),
    .C1(_05557_),
    .X(_05662_));
 sky130_fd_sc_hd__a211oi_2 _12784_ (.A1(_05599_),
    .A2(_05600_),
    .B1(_05661_),
    .C1(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__o211a_1 _12785_ (.A1(_05661_),
    .A2(_05662_),
    .B1(_05599_),
    .C1(_05600_),
    .X(_05664_));
 sky130_fd_sc_hd__o211a_1 _12786_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05559_),
    .C1(_05561_),
    .X(_05665_));
 sky130_fd_sc_hd__a211oi_2 _12787_ (.A1(_05559_),
    .A2(_05561_),
    .B1(_05663_),
    .C1(_05664_),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_1 _12788_ (.A(_05665_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _12789_ (.A(_05565_),
    .B(_05570_),
    .Y(_05668_));
 sky130_fd_sc_hd__a21oi_1 _12790_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_06427_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21a_1 _12791_ (.A1(_05667_),
    .A2(_05668_),
    .B1(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__nand3_1 _12792_ (.A(_02854_),
    .B(_02868_),
    .C(_05582_),
    .Y(_05672_));
 sky130_fd_sc_hd__a21o_1 _12793_ (.A1(_02854_),
    .A2(_05582_),
    .B1(_02868_),
    .X(_05673_));
 sky130_fd_sc_hd__a21o_1 _12794_ (.A1(_02628_),
    .A2(_05576_),
    .B1(_02596_),
    .X(_05674_));
 sky130_fd_sc_hd__nand3_1 _12795_ (.A(_02596_),
    .B(_02628_),
    .C(_05576_),
    .Y(_05675_));
 sky130_fd_sc_hd__and3_1 _12796_ (.A(_02741_),
    .B(_05674_),
    .C(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__a2bb2o_1 _12797_ (.A1_N(_05209_),
    .A2_N(_02941_),
    .B1(_02731_),
    .B2(\AuI.result[19] ),
    .X(_05677_));
 sky130_fd_sc_hd__a2bb2o_1 _12798_ (.A1_N(_02720_),
    .A2_N(_02868_),
    .B1(_03973_),
    .B2(_02742_),
    .X(_05678_));
 sky130_fd_sc_hd__a221o_1 _12799_ (.A1(\MuI.result[19] ),
    .A2(_02736_),
    .B1(_02944_),
    .B2(_05134_),
    .C1(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__a221o_1 _12800_ (.A1(\FuI.Integer[19] ),
    .A2(_04627_),
    .B1(_02718_),
    .B2(_05273_),
    .C1(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__a211o_1 _12801_ (.A1(_03110_),
    .A2(_02724_),
    .B1(_05677_),
    .C1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__a311o_1 _12802_ (.A1(_03489_),
    .A2(_05672_),
    .A3(_05673_),
    .B1(_05676_),
    .C1(_05681_),
    .X(_05683_));
 sky130_fd_sc_hd__or3_4 _12803_ (.A(_05598_),
    .B(_05670_),
    .C(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__clkbuf_1 _12804_ (.A(_05684_),
    .X(net79));
 sky130_fd_sc_hd__o21ba_1 _12805_ (.A1(_02866_),
    .A2(_05594_),
    .B1_N(_02867_),
    .X(_05685_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(_05685_),
    .A1(_02904_),
    .S(_02926_),
    .X(_05686_));
 sky130_fd_sc_hd__nand2_1 _12807_ (.A(_02805_),
    .B(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__or2_1 _12808_ (.A(_02805_),
    .B(_05686_),
    .X(_05688_));
 sky130_fd_sc_hd__and2_1 _12809_ (.A(_03271_),
    .B(_00153_),
    .X(_05689_));
 sky130_fd_sc_hd__a21oi_1 _12810_ (.A1(_03239_),
    .A2(_05959_),
    .B1(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__and3_1 _12811_ (.A(_01147_),
    .B(_05948_),
    .C(_05689_),
    .X(_05691_));
 sky130_fd_sc_hd__and4bb_1 _12812_ (.A_N(_05690_),
    .B_N(_05691_),
    .C(_00077_),
    .D(_05831_),
    .X(_05692_));
 sky130_fd_sc_hd__o2bb2a_1 _12813_ (.A1_N(_03346_),
    .A2_N(_05842_),
    .B1(_05690_),
    .B2(_05691_),
    .X(_05693_));
 sky130_fd_sc_hd__nor2_1 _12814_ (.A(_05692_),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__a21boi_1 _12815_ (.A1(_05608_),
    .A2(_05609_),
    .B1_N(_05497_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _12816_ (.A(_05617_),
    .B(_05619_),
    .Y(_05696_));
 sky130_fd_sc_hd__o2bb2a_1 _12817_ (.A1_N(_05604_),
    .A2_N(_05607_),
    .B1(_05603_),
    .B2(_05602_),
    .X(_05697_));
 sky130_fd_sc_hd__a22oi_1 _12818_ (.A1(_03443_),
    .A2(_05702_),
    .B1(_03247_),
    .B2(_00290_),
    .Y(_05698_));
 sky130_fd_sc_hd__and4_1 _12819_ (.A(_00278_),
    .B(_00279_),
    .C(_06537_),
    .D(_05756_),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_2 _12820_ (.A(_00292_),
    .B(_05649_),
    .Y(_05700_));
 sky130_fd_sc_hd__o21a_1 _12821_ (.A1(_05698_),
    .A2(_05699_),
    .B1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__nor3_1 _12822_ (.A(_05700_),
    .B(_05698_),
    .C(_05699_),
    .Y(_05703_));
 sky130_fd_sc_hd__or3_1 _12823_ (.A(_05697_),
    .B(_05701_),
    .C(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__o21ai_1 _12824_ (.A1(_05701_),
    .A2(_05703_),
    .B1(_05697_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _12825_ (.A(_05704_),
    .B(_05705_),
    .Y(_05706_));
 sky130_fd_sc_hd__xnor2_1 _12826_ (.A(_05696_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__xnor2_1 _12827_ (.A(_05695_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _12828_ (.A(_05620_),
    .B(_05622_),
    .Y(_05709_));
 sky130_fd_sc_hd__xnor2_1 _12829_ (.A(_05708_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__or2b_1 _12830_ (.A(_05624_),
    .B_N(_05626_),
    .X(_05711_));
 sky130_fd_sc_hd__xnor2_1 _12831_ (.A(_05710_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__or2b_1 _12832_ (.A(_05636_),
    .B_N(_05635_),
    .X(_05714_));
 sky130_fd_sc_hd__nand3_1 _12833_ (.A(_03733_),
    .B(_05327_),
    .C(_05637_),
    .Y(_05715_));
 sky130_fd_sc_hd__a22oi_1 _12834_ (.A1(_06442_),
    .A2(_03051_),
    .B1(_03071_),
    .B2(_06444_),
    .Y(_05716_));
 sky130_fd_sc_hd__and4_1 _12835_ (.A(_00506_),
    .B(_00676_),
    .C(_05509_),
    .D(_05574_),
    .X(_05717_));
 sky130_fd_sc_hd__nor2_1 _12836_ (.A(_05716_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__nand2_1 _12837_ (.A(_03658_),
    .B(_05456_),
    .Y(_05719_));
 sky130_fd_sc_hd__xnor2_1 _12838_ (.A(_05718_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ba_1 _12839_ (.A1(_05631_),
    .A2(_05634_),
    .B1_N(_05632_),
    .X(_05721_));
 sky130_fd_sc_hd__xnor2_1 _12840_ (.A(_05720_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _12841_ (.A(_06429_),
    .B(_05391_),
    .Y(_05723_));
 sky130_fd_sc_hd__xor2_1 _12842_ (.A(_05722_),
    .B(_05723_),
    .X(_05725_));
 sky130_fd_sc_hd__a21oi_1 _12843_ (.A1(_05714_),
    .A2(_05715_),
    .B1(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__and3_1 _12844_ (.A(_05714_),
    .B(_05715_),
    .C(_05725_),
    .X(_05727_));
 sky130_fd_sc_hd__nor2_1 _12845_ (.A(_05726_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(_03798_),
    .B(_05327_),
    .Y(_05729_));
 sky130_fd_sc_hd__xnor2_1 _12847_ (.A(_05728_),
    .B(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__xnor2_1 _12848_ (.A(_05712_),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__nor2_1 _12849_ (.A(_05629_),
    .B(_05646_),
    .Y(_05732_));
 sky130_fd_sc_hd__xnor2_1 _12850_ (.A(_05731_),
    .B(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__xnor2_1 _12851_ (.A(_05694_),
    .B(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__xnor2_1 _12852_ (.A(_05653_),
    .B(_05734_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_1 _12853_ (.A1(_05648_),
    .A2(_05651_),
    .B1(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__or3_1 _12854_ (.A(_05648_),
    .B(_05651_),
    .C(_05736_),
    .X(_05738_));
 sky130_fd_sc_hd__and2_1 _12855_ (.A(_05737_),
    .B(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__o21ai_1 _12856_ (.A1(_05655_),
    .A2(_05658_),
    .B1(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__or3_1 _12857_ (.A(_05655_),
    .B(_05658_),
    .C(_05739_),
    .X(_05741_));
 sky130_fd_sc_hd__and2_1 _12858_ (.A(_05740_),
    .B(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__and2b_1 _12859_ (.A_N(_05640_),
    .B(_05642_),
    .X(_05743_));
 sky130_fd_sc_hd__a31oi_2 _12860_ (.A1(_03842_),
    .A2(_05273_),
    .A3(_05643_),
    .B1(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__xnor2_1 _12861_ (.A(_05742_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_1 _12862_ (.A1(_05661_),
    .A2(_05663_),
    .B1(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__or3_1 _12863_ (.A(_05661_),
    .B(_05663_),
    .C(_05745_),
    .X(_05747_));
 sky130_fd_sc_hd__and2_1 _12864_ (.A(_05746_),
    .B(_05747_),
    .X(_05748_));
 sky130_fd_sc_hd__and4_1 _12865_ (.A(_05348_),
    .B(_05482_),
    .C(_05567_),
    .D(_05667_),
    .X(_05749_));
 sky130_fd_sc_hd__nor2_1 _12866_ (.A(_05565_),
    .B(_05665_),
    .Y(_05750_));
 sky130_fd_sc_hd__a311oi_2 _12867_ (.A1(_05567_),
    .A2(_05568_),
    .A3(_05667_),
    .B1(_05750_),
    .C1(_05666_),
    .Y(_05751_));
 sky130_fd_sc_hd__a21bo_1 _12868_ (.A1(_05359_),
    .A2(_05749_),
    .B1_N(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__a21oi_1 _12869_ (.A1(_05748_),
    .A2(_05752_),
    .B1(_06428_),
    .Y(_05753_));
 sky130_fd_sc_hd__o21a_1 _12870_ (.A1(_05748_),
    .A2(_05752_),
    .B1(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__or2_1 _12871_ (.A(_02630_),
    .B(_02622_),
    .X(_05755_));
 sky130_fd_sc_hd__nand2_2 _12872_ (.A(_02039_),
    .B(_05755_),
    .Y(_05757_));
 sky130_fd_sc_hd__o21a_1 _12873_ (.A1(_02039_),
    .A2(_05755_),
    .B1(_03314_),
    .X(_05758_));
 sky130_fd_sc_hd__nor2_1 _12874_ (.A(_02856_),
    .B(_02868_),
    .Y(_05759_));
 sky130_fd_sc_hd__nor2_1 _12875_ (.A(_03974_),
    .B(_03973_),
    .Y(_05760_));
 sky130_fd_sc_hd__nor2_1 _12876_ (.A(_03110_),
    .B(_05209_),
    .Y(_05761_));
 sky130_fd_sc_hd__o2bb2a_1 _12877_ (.A1_N(_05581_),
    .A2_N(_05759_),
    .B1(_05760_),
    .B2(_05761_),
    .X(_05762_));
 sky130_fd_sc_hd__a21oi_1 _12878_ (.A1(_02805_),
    .A2(_05762_),
    .B1(_02711_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21a_1 _12879_ (.A1(_02805_),
    .A2(_05762_),
    .B1(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__a2bb2o_1 _12880_ (.A1_N(_02720_),
    .A2_N(_02805_),
    .B1(_02730_),
    .B2(\AuI.result[20] ),
    .X(_05765_));
 sky130_fd_sc_hd__a221o_1 _12881_ (.A1(_05338_),
    .A2(_02718_),
    .B1(_02721_),
    .B2(_03174_),
    .C1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a2bb2o_1 _12882_ (.A1_N(_05273_),
    .A2_N(_02727_),
    .B1(_02738_),
    .B2(\MuI.result[20] ),
    .X(_05768_));
 sky130_fd_sc_hd__a311o_1 _12883_ (.A1(_03174_),
    .A2(_05273_),
    .A3(_02745_),
    .B1(_05766_),
    .C1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__a221o_1 _12884_ (.A1(\FuI.Integer[20] ),
    .A2(_06056_),
    .B1(_04642_),
    .B2(_05209_),
    .C1(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a211o_1 _12885_ (.A1(_05757_),
    .A2(_05758_),
    .B1(_05764_),
    .C1(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__a311o_4 _12886_ (.A1(_02751_),
    .A2(_05687_),
    .A3(_05688_),
    .B1(_05754_),
    .C1(_05771_),
    .X(net81));
 sky130_fd_sc_hd__a21o_1 _12887_ (.A1(_02805_),
    .A2(_05685_),
    .B1(_02802_),
    .X(_05772_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(_05772_),
    .A1(_02906_),
    .S(_04635_),
    .X(_05773_));
 sky130_fd_sc_hd__or2_1 _12889_ (.A(_02809_),
    .B(_05773_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_1 _12890_ (.A(_02809_),
    .B(_05773_),
    .Y(_05775_));
 sky130_fd_sc_hd__or2b_1 _12891_ (.A(_05744_),
    .B_N(_05742_),
    .X(_05776_));
 sky130_fd_sc_hd__or2b_1 _12892_ (.A(_05653_),
    .B_N(_05734_),
    .X(_05778_));
 sky130_fd_sc_hd__nand2_1 _12893_ (.A(_05778_),
    .B(_05737_),
    .Y(_05779_));
 sky130_fd_sc_hd__nor2_1 _12894_ (.A(_05731_),
    .B(_05732_),
    .Y(_05780_));
 sky130_fd_sc_hd__nor3_1 _12895_ (.A(_05692_),
    .B(_05693_),
    .C(_05733_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_03346_),
    .B(_05970_),
    .Y(_05782_));
 sky130_fd_sc_hd__a22o_1 _12897_ (.A1(_03346_),
    .A2(_05906_),
    .B1(_05981_),
    .B2(_03293_),
    .X(_05783_));
 sky130_fd_sc_hd__o21a_1 _12898_ (.A1(_05603_),
    .A2(_05782_),
    .B1(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__and2b_1 _12899_ (.A_N(_05710_),
    .B(_05711_),
    .X(_05785_));
 sky130_fd_sc_hd__and2_1 _12900_ (.A(_05712_),
    .B(_05730_),
    .X(_05786_));
 sky130_fd_sc_hd__a22oi_2 _12901_ (.A1(_02984_),
    .A2(_05767_),
    .B1(_03257_),
    .B2(_02983_),
    .Y(_05787_));
 sky130_fd_sc_hd__and4_1 _12902_ (.A(_00290_),
    .B(_00289_),
    .C(_03247_),
    .D(_00783_),
    .X(_05789_));
 sky130_fd_sc_hd__nor2_1 _12903_ (.A(_05787_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _12904_ (.A(_02987_),
    .B(_05713_),
    .Y(_05791_));
 sky130_fd_sc_hd__xnor2_1 _12905_ (.A(_05790_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ai_1 _12906_ (.A1(_05691_),
    .A2(_05692_),
    .B1(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__or3_1 _12907_ (.A(_05691_),
    .B(_05692_),
    .C(_05792_),
    .X(_05794_));
 sky130_fd_sc_hd__and2_1 _12908_ (.A(_05793_),
    .B(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__nor2_1 _12909_ (.A(_05699_),
    .B(_05703_),
    .Y(_05796_));
 sky130_fd_sc_hd__xor2_1 _12910_ (.A(_05795_),
    .B(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__a21boi_1 _12911_ (.A1(_05696_),
    .A2(_05705_),
    .B1_N(_05704_),
    .Y(_05798_));
 sky130_fd_sc_hd__xnor2_1 _12912_ (.A(_05797_),
    .B(_05798_),
    .Y(_05800_));
 sky130_fd_sc_hd__and2b_1 _12913_ (.A_N(_05695_),
    .B(_05707_),
    .X(_05801_));
 sky130_fd_sc_hd__a21oi_1 _12914_ (.A1(_05708_),
    .A2(_05709_),
    .B1(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__xnor2_1 _12915_ (.A(_05800_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__a22oi_1 _12916_ (.A1(_03615_),
    .A2(_05585_),
    .B1(_05660_),
    .B2(_03550_),
    .Y(_05804_));
 sky130_fd_sc_hd__and4_1 _12917_ (.A(_03550_),
    .B(_03615_),
    .C(_05585_),
    .D(_05649_),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _12918_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(_03669_),
    .B(_05520_),
    .Y(_05807_));
 sky130_fd_sc_hd__xnor2_1 _12920_ (.A(_05806_),
    .B(_05807_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ba_1 _12921_ (.A1(_05716_),
    .A2(_05719_),
    .B1_N(_05717_),
    .X(_05809_));
 sky130_fd_sc_hd__xnor2_1 _12922_ (.A(_05808_),
    .B(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand3_1 _12923_ (.A(_03744_),
    .B(_05456_),
    .C(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__a21o_1 _12924_ (.A1(_03744_),
    .A2(_05456_),
    .B1(_05810_),
    .X(_05812_));
 sky130_fd_sc_hd__nand2_1 _12925_ (.A(_05811_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__or2b_1 _12926_ (.A(_05721_),
    .B_N(_05720_),
    .X(_05814_));
 sky130_fd_sc_hd__nand3_1 _12927_ (.A(_03744_),
    .B(_05391_),
    .C(_05722_),
    .Y(_05815_));
 sky130_fd_sc_hd__nand2_1 _12928_ (.A(_05814_),
    .B(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__xnor2_1 _12929_ (.A(_05813_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _12930_ (.A(_03798_),
    .B(_05391_),
    .Y(_05818_));
 sky130_fd_sc_hd__xnor2_1 _12931_ (.A(_05817_),
    .B(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__xnor2_1 _12932_ (.A(_05803_),
    .B(_05819_),
    .Y(_05821_));
 sky130_fd_sc_hd__o21a_1 _12933_ (.A1(_05785_),
    .A2(_05786_),
    .B1(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__nor3_1 _12934_ (.A(_05785_),
    .B(_05786_),
    .C(_05821_),
    .Y(_05823_));
 sky130_fd_sc_hd__nor2_1 _12935_ (.A(_05822_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__xor2_1 _12936_ (.A(_05784_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__o21ai_1 _12937_ (.A1(_05780_),
    .A2(_05781_),
    .B1(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__or3_1 _12938_ (.A(_05780_),
    .B(_05781_),
    .C(_05825_),
    .X(_05827_));
 sky130_fd_sc_hd__and2_1 _12939_ (.A(_05826_),
    .B(_05827_),
    .X(_05828_));
 sky130_fd_sc_hd__xnor2_1 _12940_ (.A(_05779_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__a31oi_1 _12941_ (.A1(_03831_),
    .A2(_05338_),
    .A3(_05728_),
    .B1(_05726_),
    .Y(_05830_));
 sky130_fd_sc_hd__or2_1 _12942_ (.A(_05829_),
    .B(_05830_),
    .X(_05832_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_05829_),
    .B(_05830_),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _12944_ (.A(_05832_),
    .B(_05833_),
    .Y(_05834_));
 sky130_fd_sc_hd__a21o_1 _12945_ (.A1(_05740_),
    .A2(_05776_),
    .B1(_05834_),
    .X(_05835_));
 sky130_fd_sc_hd__and3_1 _12946_ (.A(_05740_),
    .B(_05776_),
    .C(_05834_),
    .X(_05836_));
 sky130_fd_sc_hd__inv_2 _12947_ (.A(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_1 _12948_ (.A(_05835_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a21boi_1 _12949_ (.A1(_05748_),
    .A2(_05752_),
    .B1_N(_05746_),
    .Y(_05839_));
 sky130_fd_sc_hd__nand2_1 _12950_ (.A(_05838_),
    .B(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21a_1 _12951_ (.A1(_05838_),
    .A2(_05839_),
    .B1(_03133_),
    .X(_05841_));
 sky130_fd_sc_hd__a21oi_2 _12952_ (.A1(_02640_),
    .A2(_05757_),
    .B1(_01962_),
    .Y(_05843_));
 sky130_fd_sc_hd__and3_1 _12953_ (.A(_01962_),
    .B(_02640_),
    .C(_05757_),
    .X(_05844_));
 sky130_fd_sc_hd__nor2_2 _12954_ (.A(_05843_),
    .B(_05844_),
    .Y(_05845_));
 sky130_fd_sc_hd__o21a_1 _12955_ (.A1(_02805_),
    .A2(_05762_),
    .B1(_04211_),
    .X(_05846_));
 sky130_fd_sc_hd__or2_1 _12956_ (.A(_02809_),
    .B(_05846_),
    .X(_05847_));
 sky130_fd_sc_hd__nand2_1 _12957_ (.A(_02809_),
    .B(_05846_),
    .Y(_05848_));
 sky130_fd_sc_hd__a21o_1 _12958_ (.A1(_05338_),
    .A2(_02745_),
    .B1(_02722_),
    .X(_05849_));
 sky130_fd_sc_hd__a2bb2o_1 _12959_ (.A1_N(_03306_),
    .A2_N(_02809_),
    .B1(_05849_),
    .B2(_03239_),
    .X(_05850_));
 sky130_fd_sc_hd__a22o_1 _12960_ (.A1(\FuI.Integer[21] ),
    .A2(_04627_),
    .B1(_02731_),
    .B2(\AuI.result[21] ),
    .X(_05851_));
 sky130_fd_sc_hd__nor2_1 _12961_ (.A(_05338_),
    .B(_02727_),
    .Y(_05852_));
 sky130_fd_sc_hd__a221o_1 _12962_ (.A1(\MuI.result[21] ),
    .A2(_02738_),
    .B1(_02945_),
    .B2(_05273_),
    .C1(_05852_),
    .X(_05854_));
 sky130_fd_sc_hd__a211o_1 _12963_ (.A1(_05402_),
    .A2(_02719_),
    .B1(_05851_),
    .C1(_05854_),
    .X(_05855_));
 sky130_fd_sc_hd__a311o_1 _12964_ (.A1(_02935_),
    .A2(_05847_),
    .A3(_05848_),
    .B1(_05850_),
    .C1(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__a221o_1 _12965_ (.A1(_05840_),
    .A2(_05841_),
    .B1(_05845_),
    .B2(_03315_),
    .C1(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__a31o_4 _12966_ (.A1(_02751_),
    .A2(_05774_),
    .A3(_05775_),
    .B1(_05857_),
    .X(net82));
 sky130_fd_sc_hd__o31ai_1 _12967_ (.A1(_02801_),
    .A2(_05273_),
    .A3(_02806_),
    .B1(_02807_),
    .Y(_05858_));
 sky130_fd_sc_hd__a31oi_2 _12968_ (.A1(_02805_),
    .A2(_02809_),
    .A3(_05685_),
    .B1(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__mux2_1 _12969_ (.A0(_05859_),
    .A1(_02907_),
    .S(_04635_),
    .X(_05860_));
 sky130_fd_sc_hd__nand2_1 _12970_ (.A(_02908_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__or2_1 _12971_ (.A(_02908_),
    .B(_05860_),
    .X(_05862_));
 sky130_fd_sc_hd__nand2_1 _12972_ (.A(_05779_),
    .B(_05828_),
    .Y(_05864_));
 sky130_fd_sc_hd__and2_1 _12973_ (.A(_05784_),
    .B(_05824_),
    .X(_05865_));
 sky130_fd_sc_hd__or2_1 _12974_ (.A(_05797_),
    .B(_05798_),
    .X(_05866_));
 sky130_fd_sc_hd__nor2_1 _12975_ (.A(_05603_),
    .B(_05782_),
    .Y(_05867_));
 sky130_fd_sc_hd__a22oi_1 _12976_ (.A1(_03454_),
    .A2(_05831_),
    .B1(_05895_),
    .B2(_03389_),
    .Y(_05868_));
 sky130_fd_sc_hd__and2_1 _12977_ (.A(_02980_),
    .B(_03444_),
    .X(_05869_));
 sky130_fd_sc_hd__and3_1 _12978_ (.A(_03389_),
    .B(_05831_),
    .C(_05869_),
    .X(_05870_));
 sky130_fd_sc_hd__nor2_1 _12979_ (.A(_05868_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__a21oi_1 _12980_ (.A1(_03497_),
    .A2(_05777_),
    .B1(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__and3_1 _12981_ (.A(_03497_),
    .B(_05777_),
    .C(_05871_),
    .X(_05873_));
 sky130_fd_sc_hd__nor2_1 _12982_ (.A(_05872_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__xnor2_1 _12983_ (.A(_05867_),
    .B(_05874_),
    .Y(_05875_));
 sky130_fd_sc_hd__a31o_1 _12984_ (.A1(_03497_),
    .A2(_05713_),
    .A3(_05790_),
    .B1(_05789_),
    .X(_05876_));
 sky130_fd_sc_hd__xor2_1 _12985_ (.A(_05875_),
    .B(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__or2b_1 _12986_ (.A(_05796_),
    .B_N(_05795_),
    .X(_05878_));
 sky130_fd_sc_hd__nand2_1 _12987_ (.A(_05793_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__xor2_1 _12988_ (.A(_05877_),
    .B(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__xnor2_1 _12989_ (.A(_05866_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__or2b_1 _12990_ (.A(_05809_),
    .B_N(_05808_),
    .X(_05882_));
 sky130_fd_sc_hd__nand2_2 _12991_ (.A(_03550_),
    .B(_03449_),
    .Y(_05883_));
 sky130_fd_sc_hd__a21boi_1 _12992_ (.A1(_03615_),
    .A2(_05660_),
    .B1_N(_05883_),
    .Y(_05885_));
 sky130_fd_sc_hd__and4_1 _12993_ (.A(_03550_),
    .B(_03615_),
    .C(_05660_),
    .D(_05713_),
    .X(_05886_));
 sky130_fd_sc_hd__nor2_1 _12994_ (.A(_05885_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand2_1 _12995_ (.A(_03669_),
    .B(_05585_),
    .Y(_05888_));
 sky130_fd_sc_hd__xnor2_1 _12996_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ba_1 _12997_ (.A1(_05804_),
    .A2(_05807_),
    .B1_N(_05805_),
    .X(_05890_));
 sky130_fd_sc_hd__xor2_1 _12998_ (.A(_05889_),
    .B(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__nand2_1 _12999_ (.A(_03733_),
    .B(_05520_),
    .Y(_05892_));
 sky130_fd_sc_hd__xnor2_1 _13000_ (.A(_05891_),
    .B(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__a21oi_1 _13001_ (.A1(_05882_),
    .A2(_05811_),
    .B1(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__and3_1 _13002_ (.A(_05882_),
    .B(_05811_),
    .C(_05893_),
    .X(_05896_));
 sky130_fd_sc_hd__nor2_1 _13003_ (.A(_05894_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _13004_ (.A(_03798_),
    .B(_05456_),
    .Y(_05898_));
 sky130_fd_sc_hd__xor2_2 _13005_ (.A(_05897_),
    .B(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__xnor2_1 _13006_ (.A(_05881_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__or2b_1 _13007_ (.A(_05803_),
    .B_N(_05819_),
    .X(_05901_));
 sky130_fd_sc_hd__o21a_1 _13008_ (.A1(_05800_),
    .A2(_05802_),
    .B1(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__xnor2_1 _13009_ (.A(_05900_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(_05782_),
    .B(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__or2_1 _13011_ (.A(_05782_),
    .B(_05903_),
    .X(_05905_));
 sky130_fd_sc_hd__and2_1 _13012_ (.A(_05904_),
    .B(_05905_),
    .X(_05907_));
 sky130_fd_sc_hd__o21ai_1 _13013_ (.A1(_05822_),
    .A2(_05865_),
    .B1(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__or3_1 _13014_ (.A(_05822_),
    .B(_05865_),
    .C(_05907_),
    .X(_05909_));
 sky130_fd_sc_hd__and2_1 _13015_ (.A(_05908_),
    .B(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__xnor2_1 _13016_ (.A(_05826_),
    .B(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__and3_1 _13017_ (.A(_05811_),
    .B(_05812_),
    .C(_05816_),
    .X(_05912_));
 sky130_fd_sc_hd__a31o_1 _13018_ (.A1(_03831_),
    .A2(_05402_),
    .A3(_05817_),
    .B1(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__xnor2_1 _13019_ (.A(_05911_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__a21o_1 _13020_ (.A1(_05864_),
    .A2(_05832_),
    .B1(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__nand3_1 _13021_ (.A(_05864_),
    .B(_05832_),
    .C(_05914_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _13022_ (.A(_05915_),
    .B(_05916_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand3_1 _13023_ (.A(_05748_),
    .B(_05835_),
    .C(_05837_),
    .Y(_05919_));
 sky130_fd_sc_hd__inv_2 _13024_ (.A(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__a21oi_1 _13025_ (.A1(_05746_),
    .A2(_05835_),
    .B1(_05836_),
    .Y(_05921_));
 sky130_fd_sc_hd__a21oi_1 _13026_ (.A1(_05752_),
    .A2(_05920_),
    .B1(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(_05918_),
    .B(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__o21a_1 _13028_ (.A1(_05918_),
    .A2(_05922_),
    .B1(_03133_),
    .X(_05924_));
 sky130_fd_sc_hd__o21ai_4 _13029_ (.A1(_02639_),
    .A2(_05843_),
    .B1(_01847_),
    .Y(_05925_));
 sky130_fd_sc_hd__o31a_2 _13030_ (.A1(_01847_),
    .A2(_02639_),
    .A3(_05843_),
    .B1(_03314_),
    .X(_05926_));
 sky130_fd_sc_hd__and2_1 _13031_ (.A(_04677_),
    .B(_05847_),
    .X(_05927_));
 sky130_fd_sc_hd__or2_1 _13032_ (.A(_02779_),
    .B(_05927_),
    .X(_05929_));
 sky130_fd_sc_hd__nand2_1 _13033_ (.A(_02779_),
    .B(_05927_),
    .Y(_05930_));
 sky130_fd_sc_hd__a2bb2o_1 _13034_ (.A1_N(_05402_),
    .A2_N(_02941_),
    .B1(_02731_),
    .B2(\AuI.result[22] ),
    .X(_05931_));
 sky130_fd_sc_hd__a32o_1 _13035_ (.A1(_03293_),
    .A2(_05402_),
    .A3(_02742_),
    .B1(_02943_),
    .B2(_05338_),
    .X(_05932_));
 sky130_fd_sc_hd__a221o_1 _13036_ (.A1(\MuI.result[22] ),
    .A2(_02737_),
    .B1(_02707_),
    .B2(_02908_),
    .C1(_05932_),
    .X(_05933_));
 sky130_fd_sc_hd__a221o_1 _13037_ (.A1(net134),
    .A2(_04627_),
    .B1(_03675_),
    .B2(_05467_),
    .C1(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__a211o_1 _13038_ (.A1(_03293_),
    .A2(_02724_),
    .B1(_05931_),
    .C1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__a31o_1 _13039_ (.A1(_03489_),
    .A2(_05929_),
    .A3(_05930_),
    .B1(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__a221o_1 _13040_ (.A1(_05923_),
    .A2(_05924_),
    .B1(_05925_),
    .B2(_05926_),
    .C1(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__a31o_4 _13041_ (.A1(_02751_),
    .A2(_05861_),
    .A3(_05862_),
    .B1(_05937_),
    .X(net83));
 sky130_fd_sc_hd__or2b_1 _13042_ (.A(_05826_),
    .B_N(_05910_),
    .X(_05938_));
 sky130_fd_sc_hd__nand2_1 _13043_ (.A(_05911_),
    .B(_05913_),
    .Y(_05939_));
 sky130_fd_sc_hd__and2b_1 _13044_ (.A_N(_05877_),
    .B(_05879_),
    .X(_05940_));
 sky130_fd_sc_hd__a21o_1 _13045_ (.A1(_03400_),
    .A2(_05981_),
    .B1(_05869_),
    .X(_05941_));
 sky130_fd_sc_hd__and3_1 _13046_ (.A(_03400_),
    .B(_05970_),
    .C(_05869_),
    .X(_05942_));
 sky130_fd_sc_hd__inv_2 _13047_ (.A(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__and4_1 _13048_ (.A(_03497_),
    .B(_05831_),
    .C(_05941_),
    .D(_05943_),
    .X(_05944_));
 sky130_fd_sc_hd__a22oi_1 _13049_ (.A1(_03497_),
    .A2(_05842_),
    .B1(_05941_),
    .B2(_05943_),
    .Y(_05945_));
 sky130_fd_sc_hd__nor2_1 _13050_ (.A(_05944_),
    .B(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_2 _13051_ (.A1(_05870_),
    .A2(_05873_),
    .B1(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__or3_1 _13052_ (.A(_05870_),
    .B(_05873_),
    .C(_05946_),
    .X(_05949_));
 sky130_fd_sc_hd__and2_1 _13053_ (.A(_05947_),
    .B(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__and2b_1 _13054_ (.A_N(_05875_),
    .B(_05876_),
    .X(_05951_));
 sky130_fd_sc_hd__a21o_1 _13055_ (.A1(_05867_),
    .A2(_05874_),
    .B1(_05951_),
    .X(_05952_));
 sky130_fd_sc_hd__xnor2_1 _13056_ (.A(_05950_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__xnor2_1 _13057_ (.A(_05940_),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__and3_1 _13058_ (.A(_03669_),
    .B(_05585_),
    .C(_05887_),
    .X(_05955_));
 sky130_fd_sc_hd__a22o_1 _13059_ (.A1(_03615_),
    .A2(_05713_),
    .B1(_05777_),
    .B2(_03550_),
    .X(_05956_));
 sky130_fd_sc_hd__o21a_1 _13060_ (.A1(_02815_),
    .A2(_05883_),
    .B1(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__nand2_1 _13061_ (.A(_03669_),
    .B(_05660_),
    .Y(_05958_));
 sky130_fd_sc_hd__xnor2_1 _13062_ (.A(_05957_),
    .B(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__o21ai_1 _13063_ (.A1(_05886_),
    .A2(_05955_),
    .B1(_05960_),
    .Y(_05961_));
 sky130_fd_sc_hd__or3_1 _13064_ (.A(_05886_),
    .B(_05955_),
    .C(_05960_),
    .X(_05962_));
 sky130_fd_sc_hd__and2_1 _13065_ (.A(_05961_),
    .B(_05962_),
    .X(_05963_));
 sky130_fd_sc_hd__nand3_1 _13066_ (.A(_03744_),
    .B(_05585_),
    .C(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__a21o_1 _13067_ (.A1(_03744_),
    .A2(_05585_),
    .B1(_05963_),
    .X(_05965_));
 sky130_fd_sc_hd__nand2_1 _13068_ (.A(_05964_),
    .B(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__or2b_1 _13069_ (.A(_05890_),
    .B_N(_05889_),
    .X(_05967_));
 sky130_fd_sc_hd__o21ai_1 _13070_ (.A1(_05891_),
    .A2(_05892_),
    .B1(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__xnor2_1 _13071_ (.A(_05966_),
    .B(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand3_1 _13072_ (.A(_03809_),
    .B(_05520_),
    .C(_05969_),
    .Y(_05971_));
 sky130_fd_sc_hd__a21o_1 _13073_ (.A1(_03809_),
    .A2(_05520_),
    .B1(_05969_),
    .X(_05972_));
 sky130_fd_sc_hd__and2_1 _13074_ (.A(_05971_),
    .B(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__and2_1 _13075_ (.A(_05954_),
    .B(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__nor2_1 _13076_ (.A(_05954_),
    .B(_05973_),
    .Y(_05975_));
 sky130_fd_sc_hd__or2_1 _13077_ (.A(_05974_),
    .B(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__or2_1 _13078_ (.A(_05866_),
    .B(_05880_),
    .X(_05977_));
 sky130_fd_sc_hd__o21ai_1 _13079_ (.A1(_05881_),
    .A2(_05899_),
    .B1(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__xnor2_1 _13080_ (.A(_05976_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21a_1 _13081_ (.A1(_05900_),
    .A2(_05902_),
    .B1(_05905_),
    .X(_05980_));
 sky130_fd_sc_hd__xnor2_1 _13082_ (.A(_05979_),
    .B(_05980_),
    .Y(_05982_));
 sky130_fd_sc_hd__xnor2_1 _13083_ (.A(_05908_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__a31o_1 _13084_ (.A1(_03831_),
    .A2(_05467_),
    .A3(_05897_),
    .B1(_05894_),
    .X(_05984_));
 sky130_fd_sc_hd__xnor2_1 _13085_ (.A(_05983_),
    .B(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__and3_1 _13086_ (.A(_05938_),
    .B(_05939_),
    .C(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__a21oi_1 _13087_ (.A1(_05938_),
    .A2(_05939_),
    .B1(_05985_),
    .Y(_05987_));
 sky130_fd_sc_hd__or2_1 _13088_ (.A(_05986_),
    .B(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__o21a_1 _13089_ (.A1(_05918_),
    .A2(_05922_),
    .B1(_05915_),
    .X(_05989_));
 sky130_fd_sc_hd__nand2_1 _13090_ (.A(_05988_),
    .B(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__o21a_1 _13091_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_03134_),
    .X(_05991_));
 sky130_fd_sc_hd__or2b_1 _13092_ (.A(_05402_),
    .B_N(_03293_),
    .X(_05993_));
 sky130_fd_sc_hd__o21ai_1 _13093_ (.A1(_02908_),
    .A2(_05859_),
    .B1(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(_05994_),
    .A1(_02909_),
    .S(_02926_),
    .X(_05995_));
 sky130_fd_sc_hd__or2_1 _13095_ (.A(_02782_),
    .B(_05995_),
    .X(_05996_));
 sky130_fd_sc_hd__a21oi_1 _13096_ (.A1(_02782_),
    .A2(_05995_),
    .B1(_02713_),
    .Y(_05997_));
 sky130_fd_sc_hd__or2b_1 _13097_ (.A(_02643_),
    .B_N(_02638_),
    .X(_05998_));
 sky130_fd_sc_hd__nand3_2 _13098_ (.A(_02632_),
    .B(_05998_),
    .C(_05925_),
    .Y(_05999_));
 sky130_fd_sc_hd__a21o_1 _13099_ (.A1(_02632_),
    .A2(_05925_),
    .B1(_05998_),
    .X(_06000_));
 sky130_fd_sc_hd__nand2_1 _13100_ (.A(_04678_),
    .B(_05929_),
    .Y(_06001_));
 sky130_fd_sc_hd__xnor2_1 _13101_ (.A(_02782_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__o22ai_1 _13102_ (.A1(_05467_),
    .A2(_02941_),
    .B1(_02782_),
    .B2(_03306_),
    .Y(_06004_));
 sky130_fd_sc_hd__a221o_1 _13103_ (.A1(\MuI.result[23] ),
    .A2(_02739_),
    .B1(_04642_),
    .B2(_05402_),
    .C1(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__a32o_1 _13104_ (.A1(_03346_),
    .A2(_05467_),
    .A3(_02744_),
    .B1(_04627_),
    .B2(\FuI.Integer[23] ),
    .X(_06006_));
 sky130_fd_sc_hd__a22o_1 _13105_ (.A1(_05531_),
    .A2(_03675_),
    .B1(_02722_),
    .B2(_03346_),
    .X(_06007_));
 sky130_fd_sc_hd__a211o_1 _13106_ (.A1(\AuI.result[23] ),
    .A2(_02732_),
    .B1(_06006_),
    .C1(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__a211o_1 _13107_ (.A1(_03489_),
    .A2(_06002_),
    .B1(_06005_),
    .C1(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__a31o_1 _13108_ (.A1(_03315_),
    .A2(_05999_),
    .A3(_06000_),
    .B1(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__a221o_4 _13109_ (.A1(_05990_),
    .A2(_05991_),
    .B1(_05996_),
    .B2(_05997_),
    .C1(_06010_),
    .X(net84));
 sky130_fd_sc_hd__o221ai_1 _13110_ (.A1(_02780_),
    .A2(_05993_),
    .B1(_02783_),
    .B2(_05859_),
    .C1(_02781_),
    .Y(_06011_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(_06011_),
    .A1(_02910_),
    .S(_04635_),
    .X(_06012_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(_02841_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__or2_1 _13113_ (.A(_02841_),
    .B(_06012_),
    .X(_06014_));
 sky130_fd_sc_hd__or2b_1 _13114_ (.A(_05966_),
    .B_N(_05968_),
    .X(_06015_));
 sky130_fd_sc_hd__and2_2 _13115_ (.A(_03626_),
    .B(_05777_),
    .X(_06016_));
 sky130_fd_sc_hd__nand2_1 _13116_ (.A(_03561_),
    .B(_05842_),
    .Y(_06017_));
 sky130_fd_sc_hd__xnor2_1 _13117_ (.A(_06016_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(_03669_),
    .B(_05713_),
    .Y(_06019_));
 sky130_fd_sc_hd__xnor2_1 _13119_ (.A(_06018_),
    .B(_06019_),
    .Y(_06020_));
 sky130_fd_sc_hd__nor2_1 _13120_ (.A(_02815_),
    .B(_05883_),
    .Y(_06021_));
 sky130_fd_sc_hd__a31o_1 _13121_ (.A1(_03669_),
    .A2(_05660_),
    .A3(_05956_),
    .B1(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _13122_ (.A(_06020_),
    .B(_06022_),
    .Y(_06024_));
 sky130_fd_sc_hd__or2_1 _13123_ (.A(_06020_),
    .B(_06022_),
    .X(_06025_));
 sky130_fd_sc_hd__nand2_1 _13124_ (.A(_06024_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_1 _13125_ (.A(_03744_),
    .B(_05660_),
    .Y(_06027_));
 sky130_fd_sc_hd__xnor2_1 _13126_ (.A(_06026_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a21o_1 _13127_ (.A1(_05961_),
    .A2(_05964_),
    .B1(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__nand3_1 _13128_ (.A(_05961_),
    .B(_05964_),
    .C(_06028_),
    .Y(_06030_));
 sky130_fd_sc_hd__and2_1 _13129_ (.A(_06029_),
    .B(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__nand3_1 _13130_ (.A(_03809_),
    .B(_05595_),
    .C(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__a21o_1 _13131_ (.A1(_03809_),
    .A2(_05595_),
    .B1(_06031_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2_1 _13132_ (.A(_06032_),
    .B(_06033_),
    .Y(_06035_));
 sky130_fd_sc_hd__a31o_1 _13133_ (.A1(_03507_),
    .A2(_05842_),
    .A3(_05941_),
    .B1(_05942_),
    .X(_06036_));
 sky130_fd_sc_hd__a22oi_1 _13134_ (.A1(_03507_),
    .A2(_05906_),
    .B1(_05981_),
    .B2(_03454_),
    .Y(_06037_));
 sky130_fd_sc_hd__a31oi_1 _13135_ (.A1(_03507_),
    .A2(_05981_),
    .A3(_05869_),
    .B1(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__and2_1 _13136_ (.A(_06036_),
    .B(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__nor2_1 _13137_ (.A(_06036_),
    .B(_06038_),
    .Y(_06040_));
 sky130_fd_sc_hd__or2_1 _13138_ (.A(_06039_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__inv_2 _13139_ (.A(_05947_),
    .Y(_06042_));
 sky130_fd_sc_hd__and2_1 _13140_ (.A(_05950_),
    .B(_05952_),
    .X(_06043_));
 sky130_fd_sc_hd__nor2_1 _13141_ (.A(_06042_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__xnor2_1 _13142_ (.A(_06041_),
    .B(_06044_),
    .Y(_06046_));
 sky130_fd_sc_hd__xor2_1 _13143_ (.A(_06035_),
    .B(_06046_),
    .X(_06047_));
 sky130_fd_sc_hd__inv_2 _13144_ (.A(_05953_),
    .Y(_06048_));
 sky130_fd_sc_hd__a21o_1 _13145_ (.A1(_05940_),
    .A2(_06048_),
    .B1(_05974_),
    .X(_06049_));
 sky130_fd_sc_hd__xor2_1 _13146_ (.A(_06047_),
    .B(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__and2b_1 _13147_ (.A_N(_05976_),
    .B(_05978_),
    .X(_06051_));
 sky130_fd_sc_hd__and2b_1 _13148_ (.A_N(_05980_),
    .B(_05979_),
    .X(_06052_));
 sky130_fd_sc_hd__or2_1 _13149_ (.A(_06051_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__xnor2_1 _13150_ (.A(_06050_),
    .B(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__a21oi_1 _13151_ (.A1(_06015_),
    .A2(_05971_),
    .B1(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__and3_1 _13152_ (.A(_06015_),
    .B(_05971_),
    .C(_06054_),
    .X(_06057_));
 sky130_fd_sc_hd__or2_1 _13153_ (.A(_06055_),
    .B(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__and2b_1 _13154_ (.A_N(_05908_),
    .B(_05982_),
    .X(_06059_));
 sky130_fd_sc_hd__a21oi_1 _13155_ (.A1(_05983_),
    .A2(_05984_),
    .B1(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nor2_2 _13156_ (.A(_06058_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__and2_1 _13157_ (.A(_06058_),
    .B(_06060_),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_1 _13158_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__or2_1 _13159_ (.A(_05918_),
    .B(_05988_),
    .X(_06064_));
 sky130_fd_sc_hd__or2_1 _13160_ (.A(_05919_),
    .B(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__or4b_1 _13161_ (.A(_05357_),
    .B(_06065_),
    .C(_05358_),
    .D_N(_05749_),
    .X(_06066_));
 sky130_fd_sc_hd__or3b_1 _13162_ (.A(_05918_),
    .B(_05988_),
    .C_N(_05921_),
    .X(_06068_));
 sky130_fd_sc_hd__o21ba_1 _13163_ (.A1(_05915_),
    .A2(_05986_),
    .B1_N(_05987_),
    .X(_06069_));
 sky130_fd_sc_hd__o311a_1 _13164_ (.A1(_05751_),
    .A2(_05919_),
    .A3(_06064_),
    .B1(_06068_),
    .C1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(_06066_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__nand2_1 _13166_ (.A(_06063_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__or2_1 _13167_ (.A(_06063_),
    .B(_06071_),
    .X(_06073_));
 sky130_fd_sc_hd__nor2_1 _13168_ (.A(_03346_),
    .B(_05467_),
    .Y(_06074_));
 sky130_fd_sc_hd__a21o_1 _13169_ (.A1(_04678_),
    .A2(_05052_),
    .B1(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__or2_1 _13170_ (.A(_02779_),
    .B(_02782_),
    .X(_06076_));
 sky130_fd_sc_hd__or4_1 _13171_ (.A(_02805_),
    .B(_02809_),
    .C(_05762_),
    .D(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__nor2_1 _13172_ (.A(_03239_),
    .B(_05338_),
    .Y(_06079_));
 sky130_fd_sc_hd__a211o_1 _13173_ (.A1(_04211_),
    .A2(_04677_),
    .B1(_06079_),
    .C1(_06076_),
    .X(_06080_));
 sky130_fd_sc_hd__nand4_1 _13174_ (.A(_02841_),
    .B(_06075_),
    .C(_06077_),
    .D(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__a31o_1 _13175_ (.A1(_06075_),
    .A2(_06077_),
    .A3(_06080_),
    .B1(_02841_),
    .X(_06082_));
 sky130_fd_sc_hd__a2bb2o_1 _13176_ (.A1_N(_05531_),
    .A2_N(_02726_),
    .B1(_02730_),
    .B2(\AuI.result[24] ),
    .X(_06083_));
 sky130_fd_sc_hd__a221o_1 _13177_ (.A1(\FuI.Integer[24] ),
    .A2(_04627_),
    .B1(_02718_),
    .B2(_05595_),
    .C1(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__a32o_1 _13178_ (.A1(_03400_),
    .A2(_05531_),
    .A3(_02743_),
    .B1(_02736_),
    .B2(\MuI.result[24] ),
    .X(_06085_));
 sky130_fd_sc_hd__nor2_1 _13179_ (.A(_02708_),
    .B(_02841_),
    .Y(_06086_));
 sky130_fd_sc_hd__o21a_1 _13180_ (.A1(_03400_),
    .A2(_05531_),
    .B1(_02721_),
    .X(_06087_));
 sky130_fd_sc_hd__a2111o_1 _13181_ (.A1(_05467_),
    .A2(_02945_),
    .B1(_06085_),
    .C1(_06086_),
    .D1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__nor2_1 _13182_ (.A(_02687_),
    .B(_02688_),
    .Y(_06089_));
 sky130_fd_sc_hd__a21oi_1 _13183_ (.A1(_02645_),
    .A2(_06089_),
    .B1(_04159_),
    .Y(_06090_));
 sky130_fd_sc_hd__o21a_1 _13184_ (.A1(_02645_),
    .A2(_06089_),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__or3_1 _13185_ (.A(_06084_),
    .B(_06088_),
    .C(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__a31o_1 _13186_ (.A1(_03489_),
    .A2(_06081_),
    .A3(_06082_),
    .B1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__a31o_1 _13187_ (.A1(_03134_),
    .A2(_06072_),
    .A3(_06073_),
    .B1(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__a31o_2 _13188_ (.A1(_02751_),
    .A2(_06013_),
    .A3(_06014_),
    .B1(_06094_),
    .X(net85));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(_02841_),
    .A2(_06011_),
    .B1(_02839_),
    .X(_06095_));
 sky130_fd_sc_hd__a21o_1 _13190_ (.A1(_02841_),
    .A2(_02910_),
    .B1(_02838_),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _13191_ (.A0(_06095_),
    .A1(_06096_),
    .S(_02925_),
    .X(_06097_));
 sky130_fd_sc_hd__a21oi_1 _13192_ (.A1(_02837_),
    .A2(_06097_),
    .B1(_02713_),
    .Y(_06099_));
 sky130_fd_sc_hd__o21a_1 _13193_ (.A1(_02837_),
    .A2(_06097_),
    .B1(_06099_),
    .X(_06100_));
 sky130_fd_sc_hd__and2_1 _13194_ (.A(_06052_),
    .B(_06050_),
    .X(_06101_));
 sky130_fd_sc_hd__o211a_1 _13195_ (.A1(_05869_),
    .A2(_06039_),
    .B1(_03507_),
    .C1(_05992_),
    .X(_06102_));
 sky130_fd_sc_hd__a21oi_1 _13196_ (.A1(_03507_),
    .A2(_05992_),
    .B1(_06039_),
    .Y(_06103_));
 sky130_fd_sc_hd__or2_1 _13197_ (.A(_06102_),
    .B(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__or3_1 _13198_ (.A(_05947_),
    .B(_06041_),
    .C(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__o21ai_1 _13199_ (.A1(_05947_),
    .A2(_06041_),
    .B1(_06104_),
    .Y(_06106_));
 sky130_fd_sc_hd__and2_1 _13200_ (.A(_06105_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__nand2_2 _13201_ (.A(_03626_),
    .B(_05906_),
    .Y(_06108_));
 sky130_fd_sc_hd__a22oi_1 _13202_ (.A1(_03626_),
    .A2(_05842_),
    .B1(_05906_),
    .B2(_03561_),
    .Y(_06109_));
 sky130_fd_sc_hd__o21ba_1 _13203_ (.A1(_06017_),
    .A2(_06108_),
    .B1_N(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__nand2_1 _13204_ (.A(_03680_),
    .B(_05777_),
    .Y(_06111_));
 sky130_fd_sc_hd__xnor2_1 _13205_ (.A(_06110_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_1 _13206_ (.A(_02815_),
    .B(_06017_),
    .Y(_06113_));
 sky130_fd_sc_hd__a31o_1 _13207_ (.A1(_03680_),
    .A2(_05713_),
    .A3(_06018_),
    .B1(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__xor2_1 _13208_ (.A(_06112_),
    .B(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__nand3_1 _13209_ (.A(_03755_),
    .B(_05713_),
    .C(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__a21o_1 _13210_ (.A1(_03755_),
    .A2(_05713_),
    .B1(_06115_),
    .X(_06117_));
 sky130_fd_sc_hd__nand2_1 _13211_ (.A(_06116_),
    .B(_06117_),
    .Y(_06118_));
 sky130_fd_sc_hd__o21ai_1 _13212_ (.A1(_06026_),
    .A2(_06027_),
    .B1(_06024_),
    .Y(_06120_));
 sky130_fd_sc_hd__xnor2_1 _13213_ (.A(_06118_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand3_1 _13214_ (.A(_03809_),
    .B(_05671_),
    .C(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__a21o_1 _13215_ (.A1(_03809_),
    .A2(_05660_),
    .B1(_06121_),
    .X(_06123_));
 sky130_fd_sc_hd__and2_1 _13216_ (.A(_06122_),
    .B(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__xor2_1 _13217_ (.A(_06107_),
    .B(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__clkinv_2 _13218_ (.A(_06041_),
    .Y(_06126_));
 sky130_fd_sc_hd__a2bb2o_1 _13219_ (.A1_N(_06035_),
    .A2_N(_06046_),
    .B1(_06126_),
    .B2(_06043_),
    .X(_06127_));
 sky130_fd_sc_hd__and2_1 _13220_ (.A(_06125_),
    .B(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__nor2_1 _13221_ (.A(_06125_),
    .B(_06127_),
    .Y(_06129_));
 sky130_fd_sc_hd__nor2_1 _13222_ (.A(_06128_),
    .B(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__and2_1 _13223_ (.A(_06051_),
    .B(_06050_),
    .X(_06131_));
 sky130_fd_sc_hd__a21o_1 _13224_ (.A1(_06047_),
    .A2(_06049_),
    .B1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__xnor2_1 _13225_ (.A(_06130_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__a21o_1 _13226_ (.A1(_06029_),
    .A2(_06032_),
    .B1(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__nand3_1 _13227_ (.A(_06029_),
    .B(_06032_),
    .C(_06133_),
    .Y(_06135_));
 sky130_fd_sc_hd__and2_1 _13228_ (.A(_06134_),
    .B(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__o21a_1 _13229_ (.A1(_06055_),
    .A2(_06101_),
    .B1(_06136_),
    .X(_06137_));
 sky130_fd_sc_hd__or3_1 _13230_ (.A(_06055_),
    .B(_06136_),
    .C(_06101_),
    .X(_06138_));
 sky130_fd_sc_hd__or2b_1 _13231_ (.A(_06137_),
    .B_N(_06138_),
    .X(_06139_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(_06063_),
    .A2(_06071_),
    .B1(_06061_),
    .Y(_06141_));
 sky130_fd_sc_hd__o21ai_1 _13233_ (.A1(_06139_),
    .A2(_06141_),
    .B1(_03133_),
    .Y(_06142_));
 sky130_fd_sc_hd__a21oi_1 _13234_ (.A1(_06139_),
    .A2(_06141_),
    .B1(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__o22ai_1 _13235_ (.A1(_05595_),
    .A2(_02941_),
    .B1(_02837_),
    .B2(_03306_),
    .Y(_06144_));
 sky130_fd_sc_hd__a221o_1 _13236_ (.A1(\MuI.result[25] ),
    .A2(_02738_),
    .B1(_04642_),
    .B2(_05531_),
    .C1(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__and2_1 _13237_ (.A(_03454_),
    .B(_05595_),
    .X(_06146_));
 sky130_fd_sc_hd__a22o_1 _13238_ (.A1(\FuI.Integer[25] ),
    .A2(_06045_),
    .B1(_02744_),
    .B2(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__a221o_1 _13239_ (.A1(_05671_),
    .A2(_02719_),
    .B1(_02722_),
    .B2(_03454_),
    .C1(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__a211o_1 _13240_ (.A1(\AuI.result[25] ),
    .A2(_02732_),
    .B1(_06145_),
    .C1(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__nand2_1 _13241_ (.A(_03400_),
    .B(_05531_),
    .Y(_06150_));
 sky130_fd_sc_hd__a21oi_1 _13242_ (.A1(_06150_),
    .A2(_06082_),
    .B1(_02837_),
    .Y(_06151_));
 sky130_fd_sc_hd__a31o_1 _13243_ (.A1(_02837_),
    .A2(_06150_),
    .A3(_06082_),
    .B1(_02711_),
    .X(_06152_));
 sky130_fd_sc_hd__a21o_1 _13244_ (.A1(_02645_),
    .A2(_06089_),
    .B1(_02687_),
    .X(_06153_));
 sky130_fd_sc_hd__xnor2_1 _13245_ (.A(_02692_),
    .B(_06153_),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_2 _13246_ (.A(_02741_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__o21a_1 _13247_ (.A1(_06151_),
    .A2(_06152_),
    .B1(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__or4b_4 _13248_ (.A(_06100_),
    .B(_06143_),
    .C(_06149_),
    .D_N(_06156_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _13249_ (.A(_06157_),
    .X(net86));
 sky130_fd_sc_hd__o21bai_1 _13250_ (.A1(_02835_),
    .A2(_06095_),
    .B1_N(_02836_),
    .Y(_06158_));
 sky130_fd_sc_hd__a21oi_1 _13251_ (.A1(_02834_),
    .A2(_06096_),
    .B1(_02836_),
    .Y(_06159_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_06158_),
    .A1(_06159_),
    .S(_04635_),
    .X(_06161_));
 sky130_fd_sc_hd__or2_1 _13253_ (.A(_02833_),
    .B(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__nand2_1 _13254_ (.A(_02833_),
    .B(_06161_),
    .Y(_06163_));
 sky130_fd_sc_hd__nand2_1 _13255_ (.A(_06130_),
    .B(_06131_),
    .Y(_06164_));
 sky130_fd_sc_hd__or2b_1 _13256_ (.A(_06118_),
    .B_N(_06120_),
    .X(_06165_));
 sky130_fd_sc_hd__nand2_1 _13257_ (.A(_06165_),
    .B(_06122_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_1 _13258_ (.A(_06112_),
    .B(_06114_),
    .Y(_06167_));
 sky130_fd_sc_hd__or3_1 _13259_ (.A(_02827_),
    .B(_02875_),
    .C(_06108_),
    .X(_06168_));
 sky130_fd_sc_hd__o21ai_1 _13260_ (.A1(_02827_),
    .A2(_02875_),
    .B1(_06108_),
    .Y(_06169_));
 sky130_fd_sc_hd__nand2_1 _13261_ (.A(_03669_),
    .B(_05842_),
    .Y(_06170_));
 sky130_fd_sc_hd__a21boi_1 _13262_ (.A1(_06168_),
    .A2(_06169_),
    .B1_N(_06170_),
    .Y(_06171_));
 sky130_fd_sc_hd__and3b_1 _13263_ (.A_N(_06170_),
    .B(_06168_),
    .C(_06169_),
    .X(_06172_));
 sky130_fd_sc_hd__nor2_1 _13264_ (.A(_06171_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__o22a_1 _13265_ (.A1(_06017_),
    .A2(_06108_),
    .B1(_06111_),
    .B2(_06109_),
    .X(_06174_));
 sky130_fd_sc_hd__xnor2_1 _13266_ (.A(_06173_),
    .B(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand3_1 _13267_ (.A(_03755_),
    .B(_05788_),
    .C(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21o_1 _13268_ (.A1(_03755_),
    .A2(_05777_),
    .B1(_06175_),
    .X(_06177_));
 sky130_fd_sc_hd__nand2_1 _13269_ (.A(_06176_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__a21oi_1 _13270_ (.A1(_06167_),
    .A2(_06116_),
    .B1(_06178_),
    .Y(_06179_));
 sky130_fd_sc_hd__and3_1 _13271_ (.A(_06167_),
    .B(_06116_),
    .C(_06178_),
    .X(_06180_));
 sky130_fd_sc_hd__nor2_1 _13272_ (.A(_06179_),
    .B(_06180_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _13273_ (.A(_03809_),
    .B(_05713_),
    .Y(_06183_));
 sky130_fd_sc_hd__xnor2_1 _13274_ (.A(_06182_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _13275_ (.A(_06102_),
    .B(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__or2_1 _13276_ (.A(_06102_),
    .B(_06184_),
    .X(_06186_));
 sky130_fd_sc_hd__a21bo_1 _13277_ (.A1(_06106_),
    .A2(_06124_),
    .B1_N(_06105_),
    .X(_06187_));
 sky130_fd_sc_hd__and3_1 _13278_ (.A(_06185_),
    .B(_06186_),
    .C(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__and2_1 _13279_ (.A(_06185_),
    .B(_06186_),
    .X(_06189_));
 sky130_fd_sc_hd__nor2_1 _13280_ (.A(_06189_),
    .B(_06187_),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_1 _13281_ (.A(_06188_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__and3_1 _13282_ (.A(_06047_),
    .B(_06049_),
    .C(_06130_),
    .X(_06192_));
 sky130_fd_sc_hd__or2_1 _13283_ (.A(_06128_),
    .B(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__xnor2_1 _13284_ (.A(_06191_),
    .B(_06193_),
    .Y(_06194_));
 sky130_fd_sc_hd__xor2_1 _13285_ (.A(_06166_),
    .B(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__a21o_1 _13286_ (.A1(_06134_),
    .A2(_06164_),
    .B1(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__and3_1 _13287_ (.A(_06134_),
    .B(_06195_),
    .C(_06164_),
    .X(_06197_));
 sky130_fd_sc_hd__inv_2 _13288_ (.A(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_1 _13289_ (.A(_06196_),
    .B(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__a2111o_1 _13290_ (.A1(_06066_),
    .A2(_06070_),
    .B1(_06139_),
    .C1(_06062_),
    .D1(_06061_),
    .X(_06200_));
 sky130_fd_sc_hd__o21ai_2 _13291_ (.A1(_06061_),
    .A2(_06137_),
    .B1(_06138_),
    .Y(_06201_));
 sky130_fd_sc_hd__nand3_1 _13292_ (.A(_06199_),
    .B(_06200_),
    .C(_06201_),
    .Y(_06203_));
 sky130_fd_sc_hd__a21o_1 _13293_ (.A1(_06200_),
    .A2(_06201_),
    .B1(_06199_),
    .X(_06204_));
 sky130_fd_sc_hd__o21ai_1 _13294_ (.A1(_06146_),
    .A2(_06151_),
    .B1(_02833_),
    .Y(_06205_));
 sky130_fd_sc_hd__o311a_1 _13295_ (.A1(_02833_),
    .A2(_06146_),
    .A3(_06151_),
    .B1(_06205_),
    .C1(_03489_),
    .X(_06206_));
 sky130_fd_sc_hd__a21o_1 _13296_ (.A1(_02645_),
    .A2(_02693_),
    .B1(_02697_),
    .X(_06207_));
 sky130_fd_sc_hd__or2_2 _13297_ (.A(_02679_),
    .B(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__nand2_2 _13298_ (.A(_02679_),
    .B(_06207_),
    .Y(_06209_));
 sky130_fd_sc_hd__a22o_1 _13299_ (.A1(_02743_),
    .A2(_02831_),
    .B1(_02944_),
    .B2(_05595_),
    .X(_06210_));
 sky130_fd_sc_hd__a21o_1 _13300_ (.A1(\MuI.result[26] ),
    .A2(_02738_),
    .B1(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__a211oi_1 _13301_ (.A1(_02705_),
    .A2(_02831_),
    .B1(_02832_),
    .C1(_02720_),
    .Y(_06212_));
 sky130_fd_sc_hd__a221o_1 _13302_ (.A1(_05724_),
    .A2(_02718_),
    .B1(_02731_),
    .B2(\AuI.result[26] ),
    .C1(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__a2bb2o_1 _13303_ (.A1_N(_05671_),
    .A2_N(_02727_),
    .B1(_04627_),
    .B2(\FuI.Integer[26] ),
    .X(_06214_));
 sky130_fd_sc_hd__or3_1 _13304_ (.A(_06211_),
    .B(_06213_),
    .C(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__a31o_1 _13305_ (.A1(_03314_),
    .A2(_06208_),
    .A3(_06209_),
    .B1(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__a311o_1 _13306_ (.A1(_03134_),
    .A2(_06203_),
    .A3(_06204_),
    .B1(_06206_),
    .C1(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__a31o_2 _13307_ (.A1(_02751_),
    .A2(_06162_),
    .A3(_06163_),
    .B1(_06217_),
    .X(net87));
 sky130_fd_sc_hd__o21a_1 _13308_ (.A1(_02833_),
    .A2(_06158_),
    .B1(_02913_),
    .X(_06218_));
 sky130_fd_sc_hd__o21ba_1 _13309_ (.A1(_02833_),
    .A2(_06159_),
    .B1_N(_02911_),
    .X(_06219_));
 sky130_fd_sc_hd__mux2_1 _13310_ (.A0(_06218_),
    .A1(_06219_),
    .S(_02926_),
    .X(_06220_));
 sky130_fd_sc_hd__or2_1 _13311_ (.A(_02830_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__nand2_1 _13312_ (.A(_02830_),
    .B(_06220_),
    .Y(_06223_));
 sky130_fd_sc_hd__or2b_1 _13313_ (.A(_06194_),
    .B_N(_06166_),
    .X(_06224_));
 sky130_fd_sc_hd__nand2_1 _13314_ (.A(_06128_),
    .B(_06191_),
    .Y(_06225_));
 sky130_fd_sc_hd__or3_1 _13315_ (.A(_06171_),
    .B(_06172_),
    .C(_06174_),
    .X(_06226_));
 sky130_fd_sc_hd__and4_1 _13316_ (.A(_03561_),
    .B(_03626_),
    .C(_05906_),
    .D(_05981_),
    .X(_06227_));
 sky130_fd_sc_hd__nand2_1 _13317_ (.A(_03680_),
    .B(_05981_),
    .Y(_06228_));
 sky130_fd_sc_hd__a22o_1 _13318_ (.A1(_03669_),
    .A2(_05906_),
    .B1(_05981_),
    .B2(_03626_),
    .X(_06229_));
 sky130_fd_sc_hd__o21a_1 _13319_ (.A1(_06108_),
    .A2(_06228_),
    .B1(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__o21a_1 _13320_ (.A1(_06227_),
    .A2(_06172_),
    .B1(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__nor3_1 _13321_ (.A(_06227_),
    .B(_06172_),
    .C(_06230_),
    .Y(_06232_));
 sky130_fd_sc_hd__nor2_1 _13322_ (.A(_06231_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__and3_1 _13323_ (.A(_03755_),
    .B(_05842_),
    .C(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__a21oi_1 _13324_ (.A1(_03755_),
    .A2(_05842_),
    .B1(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__or2_1 _13325_ (.A(_06234_),
    .B(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__a21oi_1 _13326_ (.A1(_06226_),
    .A2(_06176_),
    .B1(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__and3_1 _13327_ (.A(_06226_),
    .B(_06176_),
    .C(_06236_),
    .X(_06238_));
 sky130_fd_sc_hd__or2_1 _13328_ (.A(_06237_),
    .B(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__nand2_1 _13329_ (.A(_03820_),
    .B(_05788_),
    .Y(_06240_));
 sky130_fd_sc_hd__nor2_1 _13330_ (.A(_06239_),
    .B(_06240_),
    .Y(_06241_));
 sky130_fd_sc_hd__and2_1 _13331_ (.A(_06239_),
    .B(_06240_),
    .X(_06242_));
 sky130_fd_sc_hd__or2_1 _13332_ (.A(_06241_),
    .B(_06242_),
    .X(_06244_));
 sky130_fd_sc_hd__inv_2 _13333_ (.A(_06188_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_1 _13334_ (.A(_06185_),
    .B(_06245_),
    .Y(_06246_));
 sky130_fd_sc_hd__xnor2_1 _13335_ (.A(_06244_),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__xor2_1 _13336_ (.A(_06225_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__a31o_1 _13337_ (.A1(_03842_),
    .A2(_05724_),
    .A3(_06182_),
    .B1(_06179_),
    .X(_06249_));
 sky130_fd_sc_hd__xor2_1 _13338_ (.A(_06248_),
    .B(_06249_),
    .X(_06250_));
 sky130_fd_sc_hd__nand2_1 _13339_ (.A(_06191_),
    .B(_06192_),
    .Y(_06251_));
 sky130_fd_sc_hd__and3_1 _13340_ (.A(_06224_),
    .B(_06250_),
    .C(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__a21o_1 _13341_ (.A1(_06224_),
    .A2(_06251_),
    .B1(_06250_),
    .X(_06253_));
 sky130_fd_sc_hd__and2b_1 _13342_ (.A_N(_06252_),
    .B(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__nand2_1 _13343_ (.A(_06196_),
    .B(_06204_),
    .Y(_06255_));
 sky130_fd_sc_hd__a21oi_1 _13344_ (.A1(_06254_),
    .A2(_06255_),
    .B1(_06428_),
    .Y(_06256_));
 sky130_fd_sc_hd__o21a_1 _13345_ (.A1(_06254_),
    .A2(_06255_),
    .B1(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__a21bo_1 _13346_ (.A1(_05700_),
    .A2(_06205_),
    .B1_N(_02830_),
    .X(_06258_));
 sky130_fd_sc_hd__or3b_1 _13347_ (.A(_02831_),
    .B(_02830_),
    .C_N(_06205_),
    .X(_06259_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(_02677_),
    .B(_06209_),
    .Y(_06260_));
 sky130_fd_sc_hd__xor2_4 _13349_ (.A(_02683_),
    .B(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__a2bb2o_1 _13350_ (.A1_N(_05724_),
    .A2_N(_02941_),
    .B1(_02731_),
    .B2(\AuI.result[27] ),
    .X(_06262_));
 sky130_fd_sc_hd__a32o_1 _13351_ (.A1(_03561_),
    .A2(_05724_),
    .A3(_02742_),
    .B1(_02943_),
    .B2(_05671_),
    .X(_06263_));
 sky130_fd_sc_hd__a221o_1 _13352_ (.A1(\MuI.result[27] ),
    .A2(_02737_),
    .B1(_04011_),
    .B2(_02830_),
    .C1(_06263_),
    .X(_06265_));
 sky130_fd_sc_hd__a221o_1 _13353_ (.A1(\FuI.Integer[27] ),
    .A2(_04627_),
    .B1(_03675_),
    .B2(_05788_),
    .C1(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__a211o_1 _13354_ (.A1(_03561_),
    .A2(_02724_),
    .B1(_06262_),
    .C1(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__a21o_1 _13355_ (.A1(_03314_),
    .A2(_06261_),
    .B1(_06267_),
    .X(_06268_));
 sky130_fd_sc_hd__a31o_1 _13356_ (.A1(_04161_),
    .A2(_06258_),
    .A3(_06259_),
    .B1(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__a311o_4 _13357_ (.A1(_02751_),
    .A2(_06221_),
    .A3(_06223_),
    .B1(_06257_),
    .C1(_06269_),
    .X(net88));
 sky130_fd_sc_hd__o21a_1 _13358_ (.A1(_06196_),
    .A2(_06252_),
    .B1(_06253_),
    .X(_06270_));
 sky130_fd_sc_hd__o21a_1 _13359_ (.A1(_06197_),
    .A2(_06252_),
    .B1(_06253_),
    .X(_06271_));
 sky130_fd_sc_hd__or2b_1 _13360_ (.A(_06225_),
    .B_N(_06247_),
    .X(_06272_));
 sky130_fd_sc_hd__or2b_1 _13361_ (.A(_06248_),
    .B_N(_06249_),
    .X(_06273_));
 sky130_fd_sc_hd__nor2_1 _13362_ (.A(_06245_),
    .B(_06244_),
    .Y(_06274_));
 sky130_fd_sc_hd__inv_2 _13363_ (.A(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_1 _13364_ (.A(_06185_),
    .B(_06244_),
    .Y(_06276_));
 sky130_fd_sc_hd__and3_1 _13365_ (.A(_03680_),
    .B(_05992_),
    .C(_06108_),
    .X(_06277_));
 sky130_fd_sc_hd__xor2_1 _13366_ (.A(_02820_),
    .B(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__o21a_1 _13367_ (.A1(_06231_),
    .A2(_06234_),
    .B1(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__nor3_1 _13368_ (.A(_06231_),
    .B(_06234_),
    .C(_06278_),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_1 _13369_ (.A(_06279_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(_03831_),
    .B(_05842_),
    .Y(_06282_));
 sky130_fd_sc_hd__xor2_1 _13371_ (.A(_06281_),
    .B(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__inv_2 _13372_ (.A(_06283_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand2_1 _13373_ (.A(_06276_),
    .B(_06285_),
    .Y(_06286_));
 sky130_fd_sc_hd__or2_1 _13374_ (.A(_06276_),
    .B(_06285_),
    .X(_06287_));
 sky130_fd_sc_hd__nand2_1 _13375_ (.A(_06286_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__nor2_1 _13376_ (.A(_06275_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__and2_1 _13377_ (.A(_06275_),
    .B(_06288_),
    .X(_06290_));
 sky130_fd_sc_hd__nor2_1 _13378_ (.A(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__o21a_1 _13379_ (.A1(_06237_),
    .A2(_06241_),
    .B1(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__nor3_1 _13380_ (.A(_06237_),
    .B(_06241_),
    .C(_06291_),
    .Y(_06293_));
 sky130_fd_sc_hd__or2_1 _13381_ (.A(_06292_),
    .B(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__a21oi_1 _13382_ (.A1(_06272_),
    .A2(_06273_),
    .B1(_06294_),
    .Y(_06296_));
 sky130_fd_sc_hd__and3_1 _13383_ (.A(_06272_),
    .B(_06273_),
    .C(_06294_),
    .X(_06297_));
 sky130_fd_sc_hd__or2_1 _13384_ (.A(_06296_),
    .B(_06297_),
    .X(_06298_));
 sky130_fd_sc_hd__a311o_1 _13385_ (.A1(_06200_),
    .A2(_06201_),
    .A3(_06270_),
    .B1(_06271_),
    .C1(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__a31o_1 _13386_ (.A1(_06200_),
    .A2(_06201_),
    .A3(_06270_),
    .B1(_06271_),
    .X(_06300_));
 sky130_fd_sc_hd__a21oi_1 _13387_ (.A1(_06298_),
    .A2(_06300_),
    .B1(_06428_),
    .Y(_06301_));
 sky130_fd_sc_hd__a21bo_1 _13388_ (.A1(_05883_),
    .A2(_06258_),
    .B1_N(_02817_),
    .X(_06302_));
 sky130_fd_sc_hd__nand3b_1 _13389_ (.A_N(_02817_),
    .B(_05883_),
    .C(_06258_),
    .Y(_06303_));
 sky130_fd_sc_hd__and2_1 _13390_ (.A(_02645_),
    .B(_02694_),
    .X(_06304_));
 sky130_fd_sc_hd__o21ai_4 _13391_ (.A1(_06304_),
    .A2(_02699_),
    .B1(_01322_),
    .Y(_06305_));
 sky130_fd_sc_hd__or3_4 _13392_ (.A(_01322_),
    .B(_06304_),
    .C(_02699_),
    .X(_06306_));
 sky130_fd_sc_hd__nand2_1 _13393_ (.A(_02705_),
    .B(_06016_),
    .Y(_06307_));
 sky130_fd_sc_hd__a32o_1 _13394_ (.A1(_02707_),
    .A2(_02816_),
    .A3(_06307_),
    .B1(_02717_),
    .B2(_05853_),
    .X(_06308_));
 sky130_fd_sc_hd__nor2_1 _13395_ (.A(_05788_),
    .B(_02726_),
    .Y(_06309_));
 sky130_fd_sc_hd__a221o_1 _13396_ (.A1(\MuI.result[28] ),
    .A2(_02736_),
    .B1(_02944_),
    .B2(_05724_),
    .C1(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__a211o_1 _13397_ (.A1(\AuI.result[28] ),
    .A2(_02731_),
    .B1(_06308_),
    .C1(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__a221o_1 _13398_ (.A1(\FuI.Integer[28] ),
    .A2(_06056_),
    .B1(_02745_),
    .B2(_06016_),
    .C1(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__a31o_1 _13399_ (.A1(_03314_),
    .A2(_06305_),
    .A3(_06306_),
    .B1(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__a31o_1 _13400_ (.A1(_04161_),
    .A2(_06302_),
    .A3(_06303_),
    .B1(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__o21ba_1 _13401_ (.A1(_02829_),
    .A2(_06218_),
    .B1_N(_02828_),
    .X(_06315_));
 sky130_fd_sc_hd__mux2_1 _13402_ (.A0(_06315_),
    .A1(_02915_),
    .S(_02926_),
    .X(_06317_));
 sky130_fd_sc_hd__nand2_1 _13403_ (.A(_02817_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__o211a_1 _13404_ (.A1(_02817_),
    .A2(_06317_),
    .B1(_06318_),
    .C1(_02750_),
    .X(_06319_));
 sky130_fd_sc_hd__a211o_4 _13405_ (.A1(_06299_),
    .A2(_06301_),
    .B1(_06314_),
    .C1(_06319_),
    .X(net89));
 sky130_fd_sc_hd__o22a_1 _13406_ (.A1(_02917_),
    .A2(_02875_),
    .B1(_06108_),
    .B2(_06228_),
    .X(_06320_));
 sky130_fd_sc_hd__and3_1 _13407_ (.A(_03680_),
    .B(_05992_),
    .C(_02820_),
    .X(_06321_));
 sky130_fd_sc_hd__nor2_1 _13408_ (.A(_06320_),
    .B(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_1 _13409_ (.A(_03842_),
    .B(_05917_),
    .Y(_06323_));
 sky130_fd_sc_hd__xnor2_1 _13410_ (.A(_06322_),
    .B(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__xnor2_1 _13411_ (.A(_06286_),
    .B(_06324_),
    .Y(_06325_));
 sky130_fd_sc_hd__a31o_1 _13412_ (.A1(_03842_),
    .A2(_05853_),
    .A3(_06281_),
    .B1(_06279_),
    .X(_06326_));
 sky130_fd_sc_hd__xor2_1 _13413_ (.A(_06325_),
    .B(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__o21a_1 _13414_ (.A1(_06289_),
    .A2(_06292_),
    .B1(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__or3_1 _13415_ (.A(_06289_),
    .B(_06292_),
    .C(_06327_),
    .X(_06329_));
 sky130_fd_sc_hd__or2b_1 _13416_ (.A(_06328_),
    .B_N(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__and2b_1 _13417_ (.A_N(_06296_),
    .B(_06299_),
    .X(_06331_));
 sky130_fd_sc_hd__nand2_1 _13418_ (.A(_06330_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__o21a_1 _13419_ (.A1(_06330_),
    .A2(_06331_),
    .B1(_03133_),
    .X(_06333_));
 sky130_fd_sc_hd__nor2_1 _13420_ (.A(_02823_),
    .B(_02824_),
    .Y(_06334_));
 sky130_fd_sc_hd__or2b_1 _13421_ (.A(_05788_),
    .B_N(_03626_),
    .X(_06335_));
 sky130_fd_sc_hd__o21a_1 _13422_ (.A1(_02817_),
    .A2(_06315_),
    .B1(_06335_),
    .X(_06337_));
 sky130_fd_sc_hd__o21bai_2 _13423_ (.A1(_02817_),
    .A2(_02915_),
    .B1_N(_02919_),
    .Y(_06338_));
 sky130_fd_sc_hd__clkinv_2 _13424_ (.A(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__mux2_1 _13425_ (.A0(_06337_),
    .A1(_06339_),
    .S(_04635_),
    .X(_06340_));
 sky130_fd_sc_hd__xnor2_1 _13426_ (.A(_06334_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__a21o_1 _13427_ (.A1(_02815_),
    .A2(_06302_),
    .B1(_06334_),
    .X(_06342_));
 sky130_fd_sc_hd__or3b_1 _13428_ (.A(_06016_),
    .B(_02825_),
    .C_N(_06302_),
    .X(_06343_));
 sky130_fd_sc_hd__nand2_1 _13429_ (.A(_01320_),
    .B(_06305_),
    .Y(_06344_));
 sky130_fd_sc_hd__xor2_4 _13430_ (.A(_01327_),
    .B(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__a21o_1 _13431_ (.A1(_05853_),
    .A2(_02745_),
    .B1(_02722_),
    .X(_06346_));
 sky130_fd_sc_hd__a22o_1 _13432_ (.A1(\FuI.Integer[29] ),
    .A2(_06045_),
    .B1(_02717_),
    .B2(_05917_),
    .X(_06347_));
 sky130_fd_sc_hd__nor2_1 _13433_ (.A(_05853_),
    .B(_02726_),
    .Y(_06348_));
 sky130_fd_sc_hd__a221o_1 _13434_ (.A1(\MuI.result[29] ),
    .A2(_02736_),
    .B1(_02730_),
    .B2(\AuI.result[29] ),
    .C1(_06348_),
    .X(_06349_));
 sky130_fd_sc_hd__a211o_1 _13435_ (.A1(_04011_),
    .A2(_02825_),
    .B1(_06347_),
    .C1(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__a221o_1 _13436_ (.A1(_05788_),
    .A2(_04642_),
    .B1(_06346_),
    .B2(_03680_),
    .C1(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__a21o_1 _13437_ (.A1(_03314_),
    .A2(_06345_),
    .B1(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__a31o_1 _13438_ (.A1(_04161_),
    .A2(_06342_),
    .A3(_06343_),
    .B1(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__a221o_4 _13439_ (.A1(_06332_),
    .A2(_06333_),
    .B1(_06341_),
    .B2(_02751_),
    .C1(_06353_),
    .X(net90));
 sky130_fd_sc_hd__a31o_1 _13440_ (.A1(_03842_),
    .A2(_05917_),
    .A3(_06322_),
    .B1(_06321_),
    .X(_06354_));
 sky130_fd_sc_hd__xnor2_1 _13441_ (.A(_02812_),
    .B(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__a32o_1 _13442_ (.A1(_06276_),
    .A2(_06285_),
    .A3(_06324_),
    .B1(_06325_),
    .B2(_06326_),
    .X(_06357_));
 sky130_fd_sc_hd__xnor2_1 _13443_ (.A(_06355_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__or2_1 _13444_ (.A(_06296_),
    .B(_06328_),
    .X(_06359_));
 sky130_fd_sc_hd__inv_2 _13445_ (.A(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__a21boi_1 _13446_ (.A1(_06299_),
    .A2(_06360_),
    .B1_N(_06329_),
    .Y(_06361_));
 sky130_fd_sc_hd__nor2_1 _13447_ (.A(_06358_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__and2_1 _13448_ (.A(_06358_),
    .B(_06361_),
    .X(_06363_));
 sky130_fd_sc_hd__or2_1 _13449_ (.A(_02820_),
    .B(_02821_),
    .X(_06364_));
 sky130_fd_sc_hd__a21oi_1 _13450_ (.A1(_06170_),
    .A2(_06342_),
    .B1(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__a311o_1 _13451_ (.A1(_06364_),
    .A2(_06170_),
    .A3(_06342_),
    .B1(_06365_),
    .C1(_02711_),
    .X(_06366_));
 sky130_fd_sc_hd__a21o_1 _13452_ (.A1(_02921_),
    .A2(_06337_),
    .B1(_02824_),
    .X(_06367_));
 sky130_fd_sc_hd__a21oi_1 _13453_ (.A1(_02921_),
    .A2(_06338_),
    .B1(_02824_),
    .Y(_06368_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(_06367_),
    .A1(_06368_),
    .S(_02926_),
    .X(_06369_));
 sky130_fd_sc_hd__or2_1 _13455_ (.A(_02822_),
    .B(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__a21oi_1 _13456_ (.A1(_02822_),
    .A2(_06369_),
    .B1(_02713_),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2_1 _13457_ (.A(_01322_),
    .B(_01327_),
    .Y(_06372_));
 sky130_fd_sc_hd__nor2_1 _13458_ (.A(_06304_),
    .B(_02699_),
    .Y(_06373_));
 sky130_fd_sc_hd__o21bai_1 _13459_ (.A1(_06372_),
    .A2(_06373_),
    .B1_N(_02700_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _13460_ (.A(_01330_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__o211a_2 _13461_ (.A1(_01330_),
    .A2(_06374_),
    .B1(_06375_),
    .C1(_02741_),
    .X(_06376_));
 sky130_fd_sc_hd__a211oi_1 _13462_ (.A1(_02705_),
    .A2(_02820_),
    .B1(_02821_),
    .C1(_03306_),
    .Y(_06378_));
 sky130_fd_sc_hd__a221o_1 _13463_ (.A1(\FuI.Integer[30] ),
    .A2(_02931_),
    .B1(_02938_),
    .B2(\AuI.result[30] ),
    .C1(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__a22o_1 _13464_ (.A1(_05992_),
    .A2(_02719_),
    .B1(_04642_),
    .B2(_05853_),
    .X(_06380_));
 sky130_fd_sc_hd__nor2_1 _13465_ (.A(_05917_),
    .B(_02728_),
    .Y(_06381_));
 sky130_fd_sc_hd__a221o_1 _13466_ (.A1(\MuI.result[30] ),
    .A2(_02739_),
    .B1(_02745_),
    .B2(_02820_),
    .C1(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__or4_1 _13467_ (.A(_06376_),
    .B(_06379_),
    .C(_06380_),
    .D(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a21oi_1 _13468_ (.A1(_06370_),
    .A2(_06371_),
    .B1(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__o311ai_4 _13469_ (.A1(_06428_),
    .A2(_06362_),
    .A3(_06363_),
    .B1(_06366_),
    .C1(_06384_),
    .Y(net92));
 sky130_fd_sc_hd__o21ai_1 _13470_ (.A1(_02820_),
    .A2(_06365_),
    .B1(_02814_),
    .Y(_06385_));
 sky130_fd_sc_hd__or3_1 _13471_ (.A(_02814_),
    .B(_02820_),
    .C(_06365_),
    .X(_06386_));
 sky130_fd_sc_hd__o21ai_1 _13472_ (.A1(_02822_),
    .A2(_06367_),
    .B1(_02920_),
    .Y(_06387_));
 sky130_fd_sc_hd__a21o_1 _13473_ (.A1(_02921_),
    .A2(_06338_),
    .B1(_02824_),
    .X(_06388_));
 sky130_fd_sc_hd__a21o_1 _13474_ (.A1(_06364_),
    .A2(_06388_),
    .B1(_02918_),
    .X(_06389_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(_06387_),
    .A1(_06389_),
    .S(_04635_),
    .X(_06390_));
 sky130_fd_sc_hd__nor2_1 _13476_ (.A(_00955_),
    .B(_00956_),
    .Y(_06391_));
 sky130_fd_sc_hd__nor2_1 _13477_ (.A(_01328_),
    .B(_01329_),
    .Y(_06392_));
 sky130_fd_sc_hd__a21oi_1 _13478_ (.A1(_01330_),
    .A2(_06374_),
    .B1(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__or2_2 _13479_ (.A(_06391_),
    .B(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__nand2_2 _13480_ (.A(_06391_),
    .B(_06393_),
    .Y(_06395_));
 sky130_fd_sc_hd__a2bb2o_1 _13481_ (.A1_N(_05992_),
    .A2_N(_02728_),
    .B1(_02931_),
    .B2(\FuI.Integer[31] ),
    .X(_06396_));
 sky130_fd_sc_hd__nand2_1 _13482_ (.A(_02705_),
    .B(_02812_),
    .Y(_06398_));
 sky130_fd_sc_hd__and3_1 _13483_ (.A(_02707_),
    .B(_02813_),
    .C(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__a221o_1 _13484_ (.A1(_02744_),
    .A2(_02812_),
    .B1(_02945_),
    .B2(_05917_),
    .C1(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__a221o_1 _13485_ (.A1(\MuI.result[31] ),
    .A2(_02739_),
    .B1(_02938_),
    .B2(\AuI.result[31] ),
    .C1(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__a311o_1 _13486_ (.A1(_02741_),
    .A2(_06394_),
    .A3(_06395_),
    .B1(_06396_),
    .C1(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__a31o_1 _13487_ (.A1(_02750_),
    .A2(_02814_),
    .A3(_06390_),
    .B1(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__and2_1 _13488_ (.A(_02812_),
    .B(_06354_),
    .X(_06404_));
 sky130_fd_sc_hd__and2b_1 _13489_ (.A_N(_06355_),
    .B(_06357_),
    .X(_06405_));
 sky130_fd_sc_hd__nand3_1 _13490_ (.A(_06404_),
    .B(_06358_),
    .C(_06361_),
    .Y(_06406_));
 sky130_fd_sc_hd__o311a_1 _13491_ (.A1(_06404_),
    .A2(_06405_),
    .A3(_06363_),
    .B1(_06406_),
    .C1(_03134_),
    .X(_06407_));
 sky130_fd_sc_hd__a311o_4 _13492_ (.A1(_04161_),
    .A2(_06385_),
    .A3(_06386_),
    .B1(_06403_),
    .C1(_06407_),
    .X(net93));
 sky130_fd_sc_hd__and3_4 _13493_ (.A(\MuI.Underflow ),
    .B(_02042_),
    .C(_02151_),
    .X(_06408_));
 sky130_fd_sc_hd__clkbuf_1 _13494_ (.A(_06408_),
    .X(net103));
 sky130_fd_sc_hd__or3_1 _13495_ (.A(_02812_),
    .B(_02820_),
    .C(_06365_),
    .X(_06409_));
 sky130_fd_sc_hd__a32o_4 _13496_ (.A1(_04161_),
    .A2(_02813_),
    .A3(_06409_),
    .B1(_02739_),
    .B2(\MuI.Overflow ),
    .X(net102));
 sky130_fd_sc_hd__a22o_2 _13497_ (.A1(\MuI.Exception ),
    .A2(_02739_),
    .B1(_02732_),
    .B2(\AuI.Exception ),
    .X(net101));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(Operation[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(Operation[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(Operation[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(Operation[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(a_operand[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(a_operand[10]),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input7 (.A(a_operand[11]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(a_operand[12]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(a_operand[13]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(a_operand[14]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(a_operand[15]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(a_operand[16]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(a_operand[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input14 (.A(a_operand[18]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(a_operand[19]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(a_operand[1]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(a_operand[20]),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(a_operand[21]),
    .X(net18));
 sky130_fd_sc_hd__buf_6 input19 (.A(a_operand[22]),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input20 (.A(a_operand[23]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(a_operand[24]),
    .X(net21));
 sky130_fd_sc_hd__buf_4 input22 (.A(a_operand[25]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(a_operand[26]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(a_operand[27]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(a_operand[28]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input26 (.A(a_operand[29]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(a_operand[2]),
    .X(net27));
 sky130_fd_sc_hd__buf_6 input28 (.A(a_operand[30]),
    .X(net28));
 sky130_fd_sc_hd__buf_8 input29 (.A(a_operand[31]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(a_operand[3]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(a_operand[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(a_operand[5]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(a_operand[6]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(a_operand[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(a_operand[8]),
    .X(net35));
 sky130_fd_sc_hd__buf_4 input36 (.A(a_operand[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(b_operand[0]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(b_operand[10]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(b_operand[11]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input40 (.A(b_operand[12]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 input41 (.A(b_operand[13]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(b_operand[14]),
    .X(net42));
 sky130_fd_sc_hd__buf_4 input43 (.A(b_operand[15]),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(b_operand[16]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(b_operand[17]),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(b_operand[18]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(b_operand[19]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(b_operand[1]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(b_operand[20]),
    .X(net49));
 sky130_fd_sc_hd__buf_6 input50 (.A(b_operand[21]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(b_operand[22]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(b_operand[23]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(b_operand[24]),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(b_operand[25]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(b_operand[26]),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(b_operand[27]),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(b_operand[28]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(b_operand[29]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(b_operand[2]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input60 (.A(b_operand[30]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(b_operand[31]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(b_operand[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(b_operand[4]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 input64 (.A(b_operand[5]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(b_operand[6]),
    .X(net65));
 sky130_fd_sc_hd__buf_6 input66 (.A(b_operand[7]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(b_operand[8]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(b_operand[9]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(ALU_Output[0]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(ALU_Output[10]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ALU_Output[11]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(ALU_Output[12]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(ALU_Output[13]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(ALU_Output[14]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(ALU_Output[15]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(ALU_Output[16]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(ALU_Output[17]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(ALU_Output[18]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(ALU_Output[19]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(ALU_Output[1]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(ALU_Output[20]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(ALU_Output[21]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(ALU_Output[22]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(ALU_Output[23]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(ALU_Output[24]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(ALU_Output[25]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(ALU_Output[26]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(ALU_Output[27]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(ALU_Output[28]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(ALU_Output[29]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(ALU_Output[2]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(ALU_Output[30]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(ALU_Output[31]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(ALU_Output[3]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(ALU_Output[4]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(ALU_Output[5]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(ALU_Output[6]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(ALU_Output[7]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(ALU_Output[8]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(ALU_Output[9]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(Exception));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(Overflow));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(Underflow));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(\FuI.a_operand[24] ),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 fanout105 (.A(\FuI.a_operand[30] ),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(net67),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net65),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net64),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(net63),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net62),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(net59),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net56),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net53),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net52),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(net5),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net48),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net47),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net46),
    .X(net118));
 sky130_fd_sc_hd__buf_6 fanout119 (.A(net45),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net43),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net42),
    .X(net121));
 sky130_fd_sc_hd__buf_6 fanout122 (.A(net39),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net33),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net32),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net31),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net30),
    .X(net126));
 sky130_fd_sc_hd__buf_2 fanout127 (.A(net27),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net26),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(net25),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net24),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout131 (.A(net24),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net16),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(net12),
    .X(net133));
 sky130_fd_sc_hd__conb_1 _13037__134 (.LO(net134));
 sky130_fd_sc_hd__conb_1 \FuI._130__136  (.LO(net136));
 sky130_fd_sc_hd__conb_1 \FuI._131__137  (.LO(net137));
 sky130_fd_sc_hd__conb_1 \FuI._132__138  (.LO(net138));
 sky130_fd_sc_hd__conb_1 \FuI._133__139  (.LO(net139));
 sky130_fd_sc_hd__conb_1 \FuI._134__140  (.LO(net140));
 sky130_fd_sc_hd__conb_1 \FuI._135__141  (.LO(net141));
 sky130_fd_sc_hd__conb_1 \FuI._136__142  (.LO(net142));
 sky130_fd_sc_hd__conb_1 \FuI._137__143  (.LO(net143));
 sky130_fd_sc_hd__conb_1 \FuI._138__144  (.LO(net144));
 sky130_fd_sc_hd__conb_1 \FuI._139__145  (.LO(net145));
 sky130_fd_sc_hd__conb_1 \FuI._140__146  (.LO(net146));
 sky130_fd_sc_hd__conb_1 \FuI._141__147  (.LO(net147));
 sky130_fd_sc_hd__conb_1 \FuI._142__148  (.LO(net148));
 sky130_fd_sc_hd__conb_1 \FuI._143__149  (.LO(net149));
 sky130_fd_sc_hd__conb_1 \FuI._144__150  (.LO(net150));
 sky130_fd_sc_hd__conb_1 \FuI._145__151  (.LO(net151));
 sky130_fd_sc_hd__conb_1 \FuI._146__152  (.LO(net152));
 sky130_fd_sc_hd__conb_1 \FuI._147__153  (.LO(net153));
 sky130_fd_sc_hd__conb_1 \FuI._148__154  (.LO(net154));
 sky130_fd_sc_hd__conb_1 \FuI._149__155  (.LO(net155));
 sky130_fd_sc_hd__conb_1 \FuI._150__156  (.LO(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1607__B1_N  (.DIODE(\AuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1531__B1_N  (.DIODE(\AuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1675__C1  (.DIODE(\AuI._0024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1673__A1  (.DIODE(\AuI._0116_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1512__A  (.DIODE(\AuI._0116_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0925__A  (.DIODE(\AuI._0116_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0897__B  (.DIODE(\AuI._0116_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1675__A2  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1396__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1386__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1374__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1367__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1356__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1347__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0921__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0917__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0907__S  (.DIODE(\AuI._0126_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0908__A  (.DIODE(\AuI._0127_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0914__A  (.DIODE(\AuI._0132_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0922__A  (.DIODE(\AuI._0136_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1674__C  (.DIODE(\AuI._0138_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1043__B  (.DIODE(\AuI._0138_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0927__B  (.DIODE(\AuI._0138_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1410__A  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1354__B1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1346__B1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1275__B1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1223__C1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1209__B1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1090__A1  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1089__A  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1042__A  (.DIODE(\AuI._0139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1446__B  (.DIODE(\AuI._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1438__B  (.DIODE(\AuI._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1285__B  (.DIODE(\AuI._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1278__B  (.DIODE(\AuI._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1444__B  (.DIODE(\AuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1441__B  (.DIODE(\AuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1437__B  (.DIODE(\AuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1296__B1  (.DIODE(\AuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1295__D  (.DIODE(\AuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1494__A2  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1493__B  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1409__B  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1385__A2  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1384__B  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1364__C  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1352__A  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1327__A  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1306__A  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1303__A  (.DIODE(\AuI._0498_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1440__B  (.DIODE(\AuI._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1435__B  (.DIODE(\AuI._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1310__B1  (.DIODE(\AuI._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1309__D  (.DIODE(\AuI._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1443__A2  (.DIODE(\AuI._0519_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1439__B  (.DIODE(\AuI._0519_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1436__A2  (.DIODE(\AuI._0519_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1324__B1  (.DIODE(\AuI._0519_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1323__D  (.DIODE(\AuI._0519_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1490__B  (.DIODE(\AuI._0542_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1488__B  (.DIODE(\AuI._0542_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1349__B1  (.DIODE(\AuI._0542_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1348__C  (.DIODE(\AuI._0542_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1432__B1  (.DIODE(\AuI._0550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1428__B_N  (.DIODE(\AuI._0550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1362__B  (.DIODE(\AuI._0550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1357__B  (.DIODE(\AuI._0550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1430__A  (.DIODE(\AuI._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1429__B_N  (.DIODE(\AuI._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1427__A_N  (.DIODE(\AuI._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1369__B1  (.DIODE(\AuI._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1368__D  (.DIODE(\AuI._0560_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1503__B  (.DIODE(\AuI._0586_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1502__B  (.DIODE(\AuI._0586_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1398__B1  (.DIODE(\AuI._0586_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1397__D  (.DIODE(\AuI._0586_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1668__A2  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1663__A2  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1659__A2  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1639__A2  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1596__A  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1538__A  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1525__A  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1517__A  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1509__A  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1411__B1  (.DIODE(\AuI._0599_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._800__B1  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._799__A  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1648__B1  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1415__C  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1406__D  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0937__B_N  (.DIODE(\AuI.operand_a[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._827__A1  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._826__A1  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._822__A  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1657__B1  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1417__B  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1405__B  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0947__B_N  (.DIODE(\AuI.operand_a[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._831__C1  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._830__A  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1667__B1  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1511__B  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1418__C  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1405__D  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0955__B_N  (.DIODE(\AuI.operand_a[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._753__C_N  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._752__A1  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._722__A1  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._706__B2  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._667__A1  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._558__B2  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._475__A1  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._474__A  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._463__A  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._448__A  (.DIODE(\AuI.pe._013_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._731__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._584__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._542__B2  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._523__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._508__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._500__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._489__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._468__A1  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._467__A2  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._455__B  (.DIODE(\AuI.pe._020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._669__B1  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._571__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._557__B1  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._540__B1  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._532__B1  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._506__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._495__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._488__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._470__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._468__A2  (.DIODE(\AuI.pe._023_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._750__A  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._747__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._726__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._692__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._660__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._616__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._514__A  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._498__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._466__B1  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._462__A  (.DIODE(\AuI.pe._024_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._735__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._579__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._570__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._556__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._540__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._531__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._520__A2  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._462__B  (.DIODE(\AuI.pe._026_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._735__C1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._603__A1_N  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._579__B1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._570__B1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._540__C1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._531__B1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._520__C1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._509__A1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._490__A1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._479__A1  (.DIODE(\AuI.pe._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._740__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._571__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._558__A2  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._541__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._533__A2  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._521__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._507__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._496__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._489__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._479__B1  (.DIODE(\AuI.pe._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._673__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._608__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._581__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._572__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._541__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._532__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._521__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._507__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._496__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._489__A2  (.DIODE(\AuI.pe._050_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._769__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._713__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._583__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._553__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._535__B2  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._532__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._521__B2  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._498__A1  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._497__A  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._495__B2  (.DIODE(\AuI.pe._056_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._817__A3  (.DIODE(\AuI.pe._070_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._545__A2  (.DIODE(\AuI.pe._070_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._526__B  (.DIODE(\AuI.pe._070_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._515__A1  (.DIODE(\AuI.pe._070_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._743__A2  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._683__A2  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._674__B1  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._593__B  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._581__B1  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._572__B1  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._559__B1  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._542__A2  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._533__B1  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._523__A2  (.DIODE(\AuI.pe._079_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._768__A1  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._713__A2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._698__A2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._697__A1  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._637__B2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._626__A1  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._608__B2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._597__B2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._582__B2  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._531__A1  (.DIODE(\AuI.pe._089_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._658__D  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._588__A3  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._585__B  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._551__B  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._550__B  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._546__A1  (.DIODE(\AuI.pe._101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._792__A2  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._766__A  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._699__B2  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._655__A1  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._637__A1  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._620__D  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._599__A1  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._580__B2  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._556__A1  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._549__A  (.DIODE(\AuI.pe._105_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._816__A  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._767__B2  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._766__B  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._650__A1  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._628__A1  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._599__B2  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._595__A  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._587__A  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._579__A1  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._414__A  (.DIODE(\AuI.pe._378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._792__A1  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._765__B2  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._709__A  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._654__B2  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._638__A1  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._629__B2  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._557__B2  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._544__A  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._540__A1  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._429__A  (.DIODE(\AuI.pe._393_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._812__C  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._807__A  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._757__B2  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._650__B2  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._640__A1  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._598__A1  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._591__A  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._577__A  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._425__A1  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._404__A  (.DIODE(\AuI.pe.significand[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._810__D_N  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._808__A  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._700__B2  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._653__A1  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._605__A  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._562__A  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._422__A  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._404__B  (.DIODE(\AuI.pe.significand[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._753__A  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._752__B2  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._680__A  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._600__B2  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._485__C  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._474__C  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._469__A  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._448__B  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._409__B_N  (.DIODE(\AuI.pe.significand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._759__A1  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._753__B  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._710__A  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._521__A1  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._485__D  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._482__A  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._448__C  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._409__A  (.DIODE(\AuI.pe.significand[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._781__A2  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._681__B2  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._624__A  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._506__A1  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._504__B  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._494__A  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._445__A  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._408__B  (.DIODE(\AuI.pe.significand[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._781__A1  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._758__A1  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._504__A  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._501__A  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._444__A_N  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._408__A  (.DIODE(\AuI.pe.significand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._511__A  (.DIODE(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._510__A  (.DIODE(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._450__D_N  (.DIODE(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._443__A  (.DIODE(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._408__C  (.DIODE(\AuI.pe.significand[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._817__A1  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._680__B  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._667__A2  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._664__A_N  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._540__B2  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._530__A  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._525__A  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._450__A  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._443__B  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._408__D  (.DIODE(\AuI.pe.significand[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._754__A  (.DIODE(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._543__A  (.DIODE(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._441__A  (.DIODE(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._426__A  (.DIODE(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI.pe._407__A  (.DIODE(\AuI.pe.significand[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B2 (.DIODE(\AuI.result[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A1 (.DIODE(\AuI.result[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__B2 (.DIODE(\AuI.result[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__B2 (.DIODE(\AuI.result[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A1 (.DIODE(\AuI.result[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(\AuI.result[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A1 (.DIODE(\AuI.result[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A1 (.DIODE(\AuI.result[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11095__B2 (.DIODE(\AuI.result[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__B2 (.DIODE(\AuI.result[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B2 (.DIODE(\AuI.result[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__A1 (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6880__A  (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6857__C1  (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6846__A  (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6814__A  (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6789__A_N  (.DIODE(\MuI.Exception ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5713__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5269__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5156__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5119__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5102__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5096__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4999__A2  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4783__A2  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4667__A2  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4341__C  (.DIODE(\MuI._0017_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5269__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5156__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5119__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5102__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5096__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4828__B1  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4783__B1  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4667__B1  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4342__A  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4341__D  (.DIODE(\MuI._0018_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4463__B1  (.DIODE(\MuI._0019_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4345__A  (.DIODE(\MuI._0019_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4344__A_N  (.DIODE(\MuI._0019_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5714__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5554__C  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5513__D  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5465__D  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5411__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5354__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5320__D  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5195__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5101__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4343__B1  (.DIODE(\MuI._0020_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4440__A  (.DIODE(\MuI._0075_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4394__A  (.DIODE(\MuI._0075_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4440__B  (.DIODE(\MuI._0076_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4394__B  (.DIODE(\MuI._0076_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5758__B1  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5757__D  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5411__B2  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5354__A1  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5296__A  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5295__B2  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5142__B1  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5132__C  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5049__A1  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4403__D  (.DIODE(\MuI._0085_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5844__A2_N  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5675__A2  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5318__A  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5250__B  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5133__A2  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4957__D  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4884__C  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4709__D  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4521__C  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4405__B1  (.DIODE(\MuI._0088_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5347__B1  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5314__B  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5131__B  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4886__D  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4716__A2  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4591__B1  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4534__A2  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4523__D  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4418__D  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4417__B1  (.DIODE(\MuI._0101_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5585__B1  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5538__C  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5471__A2  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5459__B  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4907__A2  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4906__C  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4613__A2  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4605__B  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4542__B1  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4426__A  (.DIODE(\MuI._0111_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5684__B  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5612__A2  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5611__B  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5304__A2  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4726__A2  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4708__B2  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4614__A1  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4571__A1  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4544__D  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4427__A  (.DIODE(\MuI._0112_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4472__B  (.DIODE(\MuI._0154_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4465__B  (.DIODE(\MuI._0154_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4488__B_N  (.DIODE(\MuI._0166_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4476__B  (.DIODE(\MuI._0166_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5862__A2_N  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5778__A  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5694__A  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5298__A1  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5140__A  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5061__A  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5052__A  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4942__A2_N  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4850__A2_N  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4478__B  (.DIODE(\MuI._0168_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4485__C  (.DIODE(\MuI._0175_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4484__B1  (.DIODE(\MuI._0175_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4511__B  (.DIODE(\MuI._0182_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4491__B  (.DIODE(\MuI._0182_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4563__B  (.DIODE(\MuI._0208_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4514__B  (.DIODE(\MuI._0208_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5681__C  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5553__A1  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5463__B  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5229__B  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5174__B1  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5052__B  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4891__A2  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4715__D  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4600__C  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4533__D  (.DIODE(\MuI._0228_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5829__B  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5584__B  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5540__D  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5366__B  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5181__B1  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5082__B  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5079__B1  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4906__D  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4611__A  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4547__A  (.DIODE(\MuI._0244_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5748__C  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5610__B  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5578__B  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5520__A2  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5519__A2  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5291__C  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4985__C  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4978__A2  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4904__B  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4548__A  (.DIODE(\MuI._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5894__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5660__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5659__C  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5658__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5612__B1  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5434__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4734__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4732__A2  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4663__A1  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4549__A  (.DIODE(\MuI._0246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5764__B  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5682__B1  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5585__A2  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5553__B1  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5504__A2  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5367__A2  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5172__B  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4731__C  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4730__A2  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4603__B1  (.DIODE(\MuI._0305_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5580__A2  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5538__D  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5507__B  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5475__C  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5236__B  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5074__A2  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5072__A2  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4907__B1  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4613__B1  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4612__C  (.DIODE(\MuI._0315_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5748__D  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5742__B  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5580__B1  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5579__B  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5520__B1  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5292__A2_N  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5179__B  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4986__A2_N  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4908__D  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4616__A  (.DIODE(\MuI._0320_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5827__A2  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5544__A2  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5543__C1  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5434__B1  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5291__D  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5086__B  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4985__D  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4735__A  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4706__A  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4617__A  (.DIODE(\MuI._0321_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6259__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6170__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6150__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4084__B2  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3956__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3863__B2  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3862__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3793__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3783__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3453__A  (.DIODE(\MuI._0328_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6260__B2  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6169__B2  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6111__A1  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6040__A  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4304__A1  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4030__B2  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4029__A  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3543__A  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3491__A  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3454__A  (.DIODE(\MuI._0339_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6238__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4062__A  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3968__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3592__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3547__B2  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3524__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3497__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3486__A1  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3485__A  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3458__A  (.DIODE(\MuI._0350_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6342__A  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6341__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6305__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6253__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6098__A  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6097__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6028__A  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6027__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4734__B2  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3457__A  (.DIODE(\MuI._0372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5712__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5353__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5155__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5118__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5100__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5095__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4786__A2_N  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4784__D  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4671__B  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4669__D  (.DIODE(\MuI._0378_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5894__B1  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5660__B1  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5659__D  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5613__D  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5484__C1  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5221__B  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5220__A2  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4902__B  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4734__B1  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4707__A  (.DIODE(\MuI._0420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6648__A2  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6626__A2  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5887__B  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5826__B  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5635__B  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5633__A2_N  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5485__A2  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5222__A2  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4996__A2  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4708__A1  (.DIODE(\MuI._0421_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6380__B  (.DIODE(\MuI._0438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6230__B  (.DIODE(\MuI._0438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4427__B  (.DIODE(\MuI._0438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3847__B  (.DIODE(\MuI._0438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3463__A  (.DIODE(\MuI._0438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5552__B  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5540__C  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5504__B1  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5367__B1  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5362__B  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5065__B  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4974__A2_N  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4892__D  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4731__D  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4730__B1  (.DIODE(\MuI._0445_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6197__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6030__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4617__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4549__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4273__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4148__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4016__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3923__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3731__B  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3464__A  (.DIODE(\MuI._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6344__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6307__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6287__A2  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6255__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6100__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3642__A2  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3612__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3559__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3522__B  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3465__A  (.DIODE(\MuI._0460_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4708__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4663__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4571__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3621__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3520__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3508__B  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3496__B  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3486__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3484__A2  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3472__A  (.DIODE(\MuI._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6152__A1  (.DIODE(\MuI._0482_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3787__A1  (.DIODE(\MuI._0482_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3468__A  (.DIODE(\MuI._0482_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6152__A2  (.DIODE(\MuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3787__A2  (.DIODE(\MuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3468__B  (.DIODE(\MuI._0493_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6237__B  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6111__B2  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4309__C  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4170__C1  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3972__B  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3968__B2  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3967__B  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3589__A2  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3588__B  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3470__A  (.DIODE(\MuI._0515_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6386__C  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6203__C1  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6112__A2  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4026__B  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3592__B2  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3544__B  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3530__A2  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3529__B  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3524__B2  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3471__A  (.DIODE(\MuI._0526_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6241__B  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6238__B2  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3594__C  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3568__C  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3525__A2  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3504__C1  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3486__B1  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3482__A2  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3481__C  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3472__B  (.DIODE(\MuI._0537_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6155__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6117__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4343__A1  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4341__B  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4209__B2  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4208__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3942__B2  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3941__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3794__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3474__A  (.DIODE(\MuI._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6260__A1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6169__A1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6153__C1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4346__A  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4301__A1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4164__A  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4084__A1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4030__A1  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4029__B  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3475__A  (.DIODE(\MuI._0570_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6292__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6114__A1  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6039__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3966__A1  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3955__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3598__B2  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3597__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3549__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3547__A1  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3476__A  (.DIODE(\MuI._0581_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6205__A1  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3591__A1  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3545__A1  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3532__A  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3519__C  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3518__A2  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3508__A  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3498__B  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3497__B1  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3484__A1  (.DIODE(\MuI._0592_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6378__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6377__A1  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6228__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6227__A1  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6195__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4544__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4014__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3921__A1  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3727__B  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3478__A  (.DIODE(\MuI._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6342__B  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6341__A1  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6305__A1  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6098__B  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6097__A1  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6027__A1  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4902__A  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4734__A1  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3607__B  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3480__A  (.DIODE(\MuI._0625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4996__A1  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3606__A1  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3553__B  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3552__A1  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3519__B  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3518__A1  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3498__A  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3497__A2  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3482__A1  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3481__A  (.DIODE(\MuI._0636_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5939__A1  (.DIODE(\MuI._0725_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5022__B1  (.DIODE(\MuI._0725_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4994__A1  (.DIODE(\MuI._0725_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4991__A  (.DIODE(\MuI._0725_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5939__A2  (.DIODE(\MuI._0726_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4991__B  (.DIODE(\MuI._0726_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6243__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6092__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6091__A  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6020__A  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4907__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4138__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4137__A  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4006__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3721__B2  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3490__A  (.DIODE(\MuI._0735_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6298__B2  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6297__A  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6021__B2  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5894__B2  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4985__A  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3598__A1  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3597__B  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3547__A2  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3524__B1  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3491__B  (.DIODE(\MuI._0746_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6155__B  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6117__B  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4463__A1_N  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4344__C  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4209__A1  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3942__A1  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3941__B  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3874__A  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3800__B  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3493__A  (.DIODE(\MuI._0768_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6162__B2  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6160__A  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6156__A1  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6118__A1  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6047__A  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3877__B2  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3861__A  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3801__A1  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3770__A  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3494__A  (.DIODE(\MuI._0779_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6297__B  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6258__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6168__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6048__B2  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4351__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4350__B2  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4166__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4028__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3777__B2  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3495__A  (.DIODE(\MuI._0790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6298__A1  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4087__A1  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3598__A2  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3597__C  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3553__C  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3552__A2  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3548__B  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3519__D  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3518__B1  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3496__A  (.DIODE(\MuI._0801_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6373__A1_N  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6220__A1_N  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6191__C  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6090__A  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4605__A  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3916__A  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3842__A  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3722__C  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3716__C  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3502__A  (.DIODE(\MuI._0867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6300__A  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6248__A1  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6246__A1  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6245__A  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6019__A  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6018__A  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4732__A1  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4726__A1  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4135__A1_N  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3503__A  (.DIODE(\MuI._0878_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6176__B2  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6160__B  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4671__A  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4092__B2  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3940__A  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3877__A1  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3874__B  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3809__B2  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3808__A  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3515__A  (.DIODE(\MuI._1010_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6242__C  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6162__A1  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6116__A  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6047__B  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4462__A1  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4351__B  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4211__A  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3777__A1  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3770__B  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3516__A  (.DIODE(\MuI._1021_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6297__D  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6243__A2  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6154__A  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6048__A1  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4350__A1  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4037__B2  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4036__A  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3870__A1  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3799__A  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3517__A  (.DIODE(\MuI._1032_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6337__A2  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6298__B1  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6264__A1  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3607__C  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3606__A2  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3600__B  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3553__D  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3552__B1  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3522__A  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3520__A1  (.DIODE(\MuI._1043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6223__A1  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6185__B  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4731__B  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4730__A1  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4534__A1  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4264__A1  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4005__B  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3840__A1  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3720__B  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3527__A  (.DIODE(\MuI._1142_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6297__C  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6243__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6092__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6021__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6020__B  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4907__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4138__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4006__A1  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3597__D  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3528__A  (.DIODE(\MuI._1153_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6298__A2  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5894__A1  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5887__A  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5826__A  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4985__B  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3598__B1  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3549__B  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3547__B1  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3530__A1  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3529__A  (.DIODE(\MuI._1164_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6161__B  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5829__A  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4974__A1_N  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4892__C  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4592__C  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4523__C  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4519__A1_N  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3898__A  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3678__A  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3538__A  (.DIODE(\MuI._1263_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6258__B  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6212__A1  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6009__A  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5742__A  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4978__A1  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4120__A  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3896__A1  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3829__A  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3694__A1  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3539__A  (.DIODE(\MuI._1274_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6292__B  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6264__A2  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6078__A1  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5827__A1  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4253__A1  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4127__A1  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3594__B  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3592__A2  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3591__A2  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3544__A  (.DIODE(\MuI._1285_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6260__A2  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6011__B2  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5748__A  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5660__B2  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5659__A  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3995__B2  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3994__A  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3692__B2  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3592__B1  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3543__B  (.DIODE(\MuI._1318_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6638__A  (.DIODE(\MuI._1438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5636__A  (.DIODE(\MuI._1438_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6176__A1  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6174__B  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4786__A1_N  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4669__C  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4637__B2  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4467__A1  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4091__B  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3949__A  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3739__A  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3556__A  (.DIODE(\MuI._1461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6243__B1  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6242__D  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6186__A2  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6185__C  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6161__A  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6046__A  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4217__B2  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4036__B  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3772__A  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3558__A  (.DIODE(\MuI._1483_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6342__C  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6341__A2  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6301__A2  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6300__B  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4349__A  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4037__A1  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3621__A1  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3607__D  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3606__B1  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3559__A  (.DIODE(\MuI._1494_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5886__B  (.DIODE(\MuI._1662_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5836__B  (.DIODE(\MuI._1662_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5883__B  (.DIODE(\MuI._1666_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5840__B  (.DIODE(\MuI._1666_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6260__B1  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6011__A1  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5748__B  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5660__A1  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5659__B  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5222__A1  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5221__A  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3994__B  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3589__A1  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3588__A  (.DIODE(\MuI._1813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6671__A1  (.DIODE(\MuI._1836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6604__B  (.DIODE(\MuI._1836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6603__A_N  (.DIODE(\MuI._1836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5998__A  (.DIODE(\MuI._1836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6066__A  (.DIODE(\MuI._1848_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6005__B  (.DIODE(\MuI._1848_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6063__C  (.DIODE(\MuI._1908_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6060__B1  (.DIODE(\MuI._1908_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6393__A2  (.DIODE(\MuI._1975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6391__A2  (.DIODE(\MuI._1975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6121__B  (.DIODE(\MuI._1975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6500__B1  (.DIODE(\MuI._1993_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6138__A  (.DIODE(\MuI._1993_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6137__B1  (.DIODE(\MuI._1993_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6081__D  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4784__C  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4360__A  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3950__A1  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3949__B  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3756__A  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3755__B2  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3743__A  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3739__B  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3610__A  (.DIODE(\MuI._2055_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6190__A2  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6186__B1  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6185__D  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6011__A2  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6010__C  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4466__A  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4217__A1  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3880__A1  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3807__A  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3611__A  (.DIODE(\MuI._2066_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6342__D  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6341__B1  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6330__A1_N  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6306__A1  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6305__A2  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6246__A2  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6245__B  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4094__A1  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4035__A  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3612__A  (.DIODE(\MuI._2077_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5675__B1  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5346__B  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5140__B  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5133__B1  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5050__D  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4971__A2  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4884__D  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4591__A2  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4265__D  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3634__A  (.DIODE(\MuI._2319_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5257__A2  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4870__A2_N  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4259__A2_N  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4143__C  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4142__A2  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4139__D  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3847__A  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3727__D  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3725__B1  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3642__A1  (.DIODE(\MuI._2330_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5758__A2  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5354__B2  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5320__B  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5252__B1  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5142__A2  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5107__B  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5049__B2  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4956__B1  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4403__C  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3636__A  (.DIODE(\MuI._2341_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5115__A  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4959__A2_N  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4864__D  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4710__A2  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4585__B1  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4515__B  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4251__B1  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4137__C  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3720__D  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3637__A  (.DIODE(\MuI._2352_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5105__A  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4885__A2  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4710__B1  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4584__B  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4522__A2  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4399__B  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4265__C  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4264__A2  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4137__D  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3639__A  (.DIODE(\MuI._2374_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5706__B2  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4938__A  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4643__A  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4494__A  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4493__B2  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4373__B  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4372__A1  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3831__B1  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3830__C  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3646__C  (.DIODE(\MuI._2440_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5792__A  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5706__A1  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4850__A1_N  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4750__C  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4494__C  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4493__A2  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3913__C  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3675__C  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3653__A  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3646__D  (.DIODE(\MuI._2451_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6154__B  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6080__A  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4888__A1_N  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4717__C  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4713__A1_N  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4588__A1_N  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4399__A  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4246__A  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3993__A  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3650__A  (.DIODE(\MuI._2473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5709__A  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5263__A1  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5149__B2  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4942__A1_N  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4848__C  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4624__B1  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3838__C  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3689__A  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3675__D  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3649__A  (.DIODE(\MuI._2484_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6787__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6715__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6712__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6706__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6703__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6688__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6676__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6670__S  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6587__B  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6585__A  (.DIODE(\MuI._2486_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6776__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6747__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6743__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6737__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6736__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6731__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6725__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6721__S  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6588__A2  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6586__B1  (.DIODE(\MuI._2487_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4492__B  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4397__C  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4396__A2  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4244__D  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3914__B1  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3913__D  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3840__A2  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3688__C  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3679__B1  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3650__B  (.DIODE(\MuI._2495_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4226__A  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4118__C  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4117__A2  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4006__A2  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4005__C  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3898__B  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3704__D  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3701__B1  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3658__A  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3655__A2  (.DIODE(\MuI._2528_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6635__C  (.DIODE(\MuI._2534_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6259__C  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6162__A2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6156__A2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6010__A  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4716__B2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4251__B2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4125__B2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3688__A  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3679__B2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3655__B2  (.DIODE(\MuI._2550_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6786__B1  (.DIODE(\MuI._2559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6659__B1  (.DIODE(\MuI._2559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6787__A0  (.DIODE(\MuI._2563_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6786__A2  (.DIODE(\MuI._2563_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6659__C1  (.DIODE(\MuI._2563_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6658__D  (.DIODE(\MuI._2566_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6153__D1  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6046__B  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5684__A  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5236__A  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5179__A  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4963__A1_N  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4870__A1_N  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4116__A  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4035__B  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3671__A1  (.DIODE(\MuI._2583_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5714__A1  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4998__A  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4939__B2  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4836__A1  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4480__B  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4479__A1  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4100__B  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4099__A1  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3901__A2  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3660__A  (.DIODE(\MuI._2605_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6222__D  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4741__A  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4358__A  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4228__A  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4227__B2  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4102__A  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3899__C  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3883__B  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3670__B  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3661__A  (.DIODE(\MuI._2616_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6715__A0  (.DIODE(\MuI._2625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6712__A1  (.DIODE(\MuI._2625_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6721__A0  (.DIODE(\MuI._2629_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6715__A1  (.DIODE(\MuI._2629_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6148__C  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6117__D  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5765__B  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5237__B  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4970__B  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4884__B  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4709__B  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3949__D  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3703__A  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3663__A  (.DIODE(\MuI._2638_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5794__A  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5793__B2  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5712__A  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5157__B2  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4939__A1  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4749__B2  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4373__A  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4228__B  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3901__B1  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3665__A  (.DIODE(\MuI._2660_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4835__A  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4478__A  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4372__B2  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4227__A1  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4098__A  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3899__D  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3831__A2  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3704__C  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3670__D  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3666__A  (.DIODE(\MuI._2671_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6148__B  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6117__C  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5765__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5237__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4970__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4709__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3950__A2  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3949__C  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3702__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3668__A  (.DIODE(\MuI._2693_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6857__B1  (.DIODE(\MuI._2731_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6814__B  (.DIODE(\MuI._2731_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6810__A  (.DIODE(\MuI._2731_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6857__A2  (.DIODE(\MuI._2733_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6846__B  (.DIODE(\MuI._2733_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6814__C  (.DIODE(\MuI._2733_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6810__B_N  (.DIODE(\MuI._2733_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5265__A  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4763__A2_N  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4516__A2  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4397__D  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4125__A2  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3838__D  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3715__A2  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3712__C  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3688__D  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3678__B  (.DIODE(\MuI._2773_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4585__A2  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4516__B1  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4395__B  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4251__A2  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4125__B1  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3721__A2  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3720__C  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3715__B1  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3712__D  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3687__A  (.DIODE(\MuI._2786_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6380__A  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6098__D  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6097__B1  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6028__C  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6027__A2  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6018__B  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4243__B1  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4116__B  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4008__B  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3692__A2  (.DIODE(\MuI._2789_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5862__A1_N  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5695__A  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5195__B2  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5112__B2  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4947__C  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4760__B1  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4625__D  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4517__C  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4124__C  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3691__A  (.DIODE(\MuI._2790_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6100__A  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6028__D  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6027__B1  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4396__B1  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4242__B  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4014__C  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4012__A2  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3916__B  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3840__B1  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3692__B1  (.DIODE(\MuI._2791_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6168__B  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5848__A1_N  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5764__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4886__C  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4584__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4395__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4242__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3948__B  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3760__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3698__A  (.DIODE(\MuI._2796_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6378__D  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6377__B1  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6230__A  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6098__C  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6097__A2  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6019__B  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4006__B1  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3896__A2  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3829__B  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3698__B  (.DIODE(\MuI._2797_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5681__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5238__B2  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5180__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5046__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4971__B2  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4884__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4586__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4517__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3884__C  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3700__A  (.DIODE(\MuI._2799_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6238__B1  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6169__A2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6048__A2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5074__B2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4396__B2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4243__B2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4117__B2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4037__A2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4036__C  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3701__B2  (.DIODE(\MuI._2800_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6170__C  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6150__B  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6118__A2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5766__B2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5181__B2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4885__B2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4710__B2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4585__B2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3885__A2  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3704__A  (.DIODE(\MuI._2802_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6170__D  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6118__B1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5766__A1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5181__A1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4885__A1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4710__A1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4585__A1  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4244__B  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4118__B  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3704__B  (.DIODE(\MuI._2803_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6242__B  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6190__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6186__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6091__B  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4906__B  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4417__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4137__B  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3914__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3721__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3715__A1  (.DIODE(\MuI._2813_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6242__A  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6223__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6190__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6186__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4906__A  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4417__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4005__A  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3914__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3720__A  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3715__B2  (.DIODE(\MuI._2814_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6184__A  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4986__A1_N  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4908__C  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4904__A  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4536__A  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4259__A1_N  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4139__C  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4008__A  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3912__A  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3718__A1_N  (.DIODE(\MuI._2817_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6378__A  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6377__B2  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6228__A  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6227__B2  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4613__B2  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4612__A  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4544__A  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4421__B2  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3921__B2  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3727__A  (.DIODE(\MuI._2826_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5766__A2  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5765__C  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5673__B  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5404__A2  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5346__D  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4971__B1  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4715__C  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4590__D  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4533__C  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3730__A  (.DIODE(\MuI._2829_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5297__A2  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5058__C  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4963__A2_N  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4588__A2_N  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4269__C  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4268__A2  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4261__B  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4143__D  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4142__B1  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3731__A  (.DIODE(\MuI._2830_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5757__A  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5078__A  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5070__B2  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5067__B2  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4863__B2  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4760__B2  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4100__C  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3942__A2  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3808__C  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3739__C  (.DIODE(\MuI._2836_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5231__A1  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5230__B  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4956__A1  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4955__B  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4862__B  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4759__B  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4623__C  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3756__D  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3745__A  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3738__A  (.DIODE(\MuI._2837_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5757__B  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5174__A1  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5078__B  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5070__A1  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5067__A1  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4863__A1  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3876__A  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3874__D  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3808__D  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3739__D  (.DIODE(\MuI._2838_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6222__C  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6189__D  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4636__A  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4359__A1  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4100__A  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4099__B2  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3885__A1  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3884__B  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3816__A  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3742__A  (.DIODE(\MuI._2840_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5229__A  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5172__A  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5065__A  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4959__A1_N  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4866__A1_N  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4864__C  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4763__A1_N  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4098__B  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3873__B  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3742__B  (.DIODE(\MuI._2841_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6189__C  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6175__B  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6082__B1  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4831__A1_N  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4359__B2  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4218__B  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4213__A  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3885__B2  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3884__A  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3746__A1  (.DIODE(\MuI._2843_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5675__B2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5174__B2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5079__B2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4494__B  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4373__C  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4228__C  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4099__A2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3874__C  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3809__A2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3746__A2  (.DIODE(\MuI._2844_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5675__A1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5079__A1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4494__D  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4493__B1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4373__D  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4228__D  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4099__B1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3942__B1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3809__B1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3746__B1  (.DIODE(\MuI._2845_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6307__A  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6287__B2  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6254__A1  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6253__B1  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6220__A2_N  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6195__C  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6194__A2  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6078__A2  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6009__B  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3757__A1  (.DIODE(\MuI._2849_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5082__A  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5080__C  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5072__A1  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4492__A  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4371__A  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4226__B  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4102__B  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3880__A2  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3807__B  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3751__A  (.DIODE(\MuI._2850_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6386__B  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6203__B1  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6114__A2  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6112__A1  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6111__A2  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6039__B  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5678__A1  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5292__A1_N  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4028__B  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3757__A2  (.DIODE(\MuI._2851_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5714__B2  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5713__A  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4837__A  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4836__B2  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4742__A1  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4480__A  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4479__B2  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4360__B  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3756__B  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3755__A1  (.DIODE(\MuI._2852_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5758__B2  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5674__A  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5173__A  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5071__A  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5066__A  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4956__B2  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4624__B2  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3941__C  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3875__A  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3755__A2  (.DIODE(\MuI._2853_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5758__A1  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5674__B  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5173__B  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5071__B  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5066__B  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4760__A1  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4624__A2  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4100__D  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3941__D  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3755__B1  (.DIODE(\MuI._2854_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6241__A  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6238__A2  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6237__A  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6205__A2  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5658__A1  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5220__A1  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3992__A2  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3828__A1  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3815__A  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3761__A  (.DIODE(\MuI._2860_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5779__C  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5141__A  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5060__B2  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4945__C  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4846__C  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4748__C  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4645__C  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4644__A2  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3773__A  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3767__A  (.DIODE(\MuI._2866_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5695__B  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5423__B2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5368__A  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5367__B2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5133__B2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4359__A2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4092__A2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3863__A2  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3800__C  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3770__C  (.DIODE(\MuI._2867_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5779__D  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5141__B  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5060__A1  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4945__D  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4846__D  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4748__D  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4644__B1  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4480__D  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3775__A  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3769__A  (.DIODE(\MuI._2868_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5423__A1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5368__B  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5367__A1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5133__A1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4359__B1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4092__B1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3863__B1  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3862__D  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3800__D  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3770__D  (.DIODE(\MuI._2869_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5422__A  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5366__A  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5362__A  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5257__A1  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5131__A  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4358__B  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4213__B  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3861__B  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3798__A  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3772__B  (.DIODE(\MuI._2871_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5696__A1  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5424__A  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5251__A  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5142__B2  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5132__A  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5059__A  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5054__B2  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4479__A2  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4360__C  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3774__A  (.DIODE(\MuI._2873_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5520__B2  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5475__A  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5058__A  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4218__C  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4217__A2  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3968__B1  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3956__B  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3862__C  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3801__A2  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3777__A2  (.DIODE(\MuI._2874_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5780__B1  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5696__B1  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5695__D  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5424__B  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5251__C  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5142__A1  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5054__A1  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4479__B1  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4360__D  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3776__A  (.DIODE(\MuI._2875_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5544__A1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5543__B1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5520__A1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5475__B  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5058__B  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4218__D  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4217__B1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3957__B1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3801__B1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3777__B1  (.DIODE(\MuI._2876_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5793__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5456__A1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5403__B  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5295__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5263__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5149__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5049__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4836__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4467__B1  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3782__A  (.DIODE(\MuI._2881_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5707__C  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5295__A1  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5263__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5149__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5112__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5107__C  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5106__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4467__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4209__A2  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3786__A  (.DIODE(\MuI._2885_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6151__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6041__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4298__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3957__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3868__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3791__A2  (.DIODE(\MuI._2889_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6151__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6041__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4298__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3957__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3868__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3791__A3  (.DIODE(\MuI._2890_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5706__A2  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5539__B2  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5505__A  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5456__B2  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5404__B2  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5403__A  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5347__B2  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5346__A  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4086__C  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3793__B  (.DIODE(\MuI._2892_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6259__B  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6170__B  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6156__B2  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6118__B2  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4086__B  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3863__A1  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3862__B  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3801__B2  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3800__A  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3796__A  (.DIODE(\MuI._2894_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5459__A  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5406__A  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5349__A  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5314__A  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5199__A1_N  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5105__B  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4835__B  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4466__B  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4211__B  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3796__B  (.DIODE(\MuI._2895_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5304__A1  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4216__B  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4094__A2  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4026__A  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3968__A2  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3967__A  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3966__A2  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3955__B  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3870__A2  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3799__B  (.DIODE(\MuI._2898_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6287__A1  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6255__A  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6227__A2  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6195__D  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6194__B1  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6092__B1  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6021__A2  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3896__B2  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3828__A2  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3815__B  (.DIODE(\MuI._2914_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5681__B  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5238__A1  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5180__B  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5046__B  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4971__A1  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4586__B  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4517__B  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3950__B1  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3884__D  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3819__A  (.DIODE(\MuI._2918_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6169__B1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6048__B1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5086__A  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5074__A1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4396__A1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4243__A1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4117__A1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4037__B1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4036__D  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3820__B1  (.DIODE(\MuI._2919_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3854__A  (.DIODE(\MuI._2926_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3853__A  (.DIODE(\MuI._2926_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6189__A  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6185__A  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4731__A  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4730__B2  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4603__B2  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4534__B2  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4418__A  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4264__B2  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3913__A  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3840__B2  (.DIODE(\MuI._2939_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5792__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5709__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5541__A  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5265__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5115__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5050__C  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4938__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4741__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4636__B  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3867__A  (.DIODE(\MuI._2966_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5519__A1  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5507__A  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5471__A1  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5297__A1  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4349__B  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4166__B  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4087__A2  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4062__B  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3972__A  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3868__C1  (.DIODE(\MuI._2967_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6111__B1  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6040__B  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5434__B2  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5291__A  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4493__A1  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4372__A2  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4227__A2  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4030__A2  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4029__C  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3877__A2  (.DIODE(\MuI._2975_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6041__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5485__A1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5484__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5434__A1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5291__B  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4372__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4227__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4030__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4029__D  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3877__B1  (.DIODE(\MuI._2976_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6344__A  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6305__B1  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6253__A2  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6252__C  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6248__A2  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6212__A2  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6184__B  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6080__B  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4216__A  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3992__A1  (.DIODE(\MuI._3091_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6063__A  (.DIODE(\MuI._3154_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6060__A1  (.DIODE(\MuI._3154_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4056__A  (.DIODE(\MuI._3154_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5999__B  (.DIODE(\MuI._3156_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4057__B  (.DIODE(\MuI._3156_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4078__B  (.DIODE(\MuI._3158_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4076__A  (.DIODE(\MuI._3158_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4183__A  (.DIODE(\MuI._3160_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4074__A  (.DIODE(\MuI._3160_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4072__A  (.DIODE(\MuI._3160_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4183__B  (.DIODE(\MuI._3171_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4074__B  (.DIODE(\MuI._3171_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4072__B  (.DIODE(\MuI._3171_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5706__B1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5539__A1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5505__B  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5404__A1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5347__A2  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5346__C  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5112__B1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5106__B1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4209__B1  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4086__D  (.DIODE(\MuI._3185_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5780__A2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5303__A  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5302__B2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5252__B2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5053__A  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4946__A2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4847__A2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4749__A2  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4480__C  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4091__C  (.DIODE(\MuI._3189_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5303__B  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5302__A1  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5252__A2  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5132__B  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5059__B  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5053__B  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4946__B1  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4847__B1  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4749__B1  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4091__D  (.DIODE(\MuI._3190_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5778__B  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5695__C  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5152__A  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5106__B2  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4866__A2_N  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4761__D  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4586__C  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4517__D  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4250__C  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4124__D  (.DIODE(\MuI._3223_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5766__B1  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5682__A2  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5404__B1  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5349__B  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4972__D  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4716__B1  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4603__A2  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4592__D  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4534__B1  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4147__A  (.DIODE(\MuI._3246_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5848__A2_N  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5678__A2  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5058__D  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4713__A2_N  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4422__C  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4421__A2  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4414__B  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4269__D  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4268__B1  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4148__A  (.DIODE(\MuI._3247_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5714__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5513__B  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5465__C  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5464__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5411__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5354__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5320__C  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5319__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5195__A2  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4163__B  (.DIODE(\MuI._3262_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5552__A  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5511__A  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5463__A  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5410__B  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5318__B  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5194__B  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4831__A2_N  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4463__A2_N  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4344__D  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4169__A  (.DIODE(\MuI._3268_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5633__A1_N  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5613__C  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5584__A  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4462__A2  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4346__B  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4309__B  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4305__A1  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4304__A2  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4301__A2  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4170__B1  (.DIODE(\MuI._3269_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4181__A  (.DIODE(\MuI._3278_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4180__A  (.DIODE(\MuI._3278_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4181__B  (.DIODE(\MuI._3279_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4180__B  (.DIODE(\MuI._3279_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5794__C  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5793__A2  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5457__A  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5296__B  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5262__C  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5150__C  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5113__C  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5049__A2  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4836__A2  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4208__C  (.DIODE(\MuI._3306_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5707__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5457__B  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5296__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5262__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5150__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5113__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5107__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4939__B1  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4637__B1  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4208__D  (.DIODE(\MuI._3307_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5757__C  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5694__B  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5319__A1  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5251__D  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5194__A  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5106__A1  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4709__C  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4586__D  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4405__A2  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4250__D  (.DIODE(\MuI._3349_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5756__B  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5464__B2  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5411__A1  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5353__A  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5295__A2  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5054__A2  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4970__C  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4590__C  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4521__D  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4263__A  (.DIODE(\MuI._3362_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5347__A1  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5199__A2_N  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4885__B1  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4711__D  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4522__B1  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4519__A2_N  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4418__C  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4417__A2  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4406__D  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4264__B1  (.DIODE(\MuI._3363_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5681__D  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5586__C  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5511__B  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5505__C  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5368__C  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5298__A2  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5061__B  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4891__B1  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4600__D  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4272__A  (.DIODE(\MuI._3371_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5406__B  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4888__A2_N  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4717__D  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4606__B  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4544__C  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4542__A2  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4536__B  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4422__D  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4421__B1  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4273__A  (.DIODE(\MuI._3372_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5713__D  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5412__D  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5355__D  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5270__B1  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5196__D  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5157__B1  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5120__B1  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5097__B1  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4999__B1  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4297__A  (.DIODE(\MuI._3396_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6626__A1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5612__A1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5610__A  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5586__B  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5585__A1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5553__A2  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5512__B1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5464__B1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5319__B1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4298__B1  (.DIODE(\MuI._3397_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5412__C  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5355__C  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5270__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5196__C  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5157__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5120__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5101__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5097__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4343__A2  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4303__A  (.DIODE(\MuI._3402_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4322__A_N  (.DIODE(\MuI._3418_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4321__A  (.DIODE(\MuI._3418_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4322__B  (.DIODE(\MuI._3420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4321__B  (.DIODE(\MuI._3420_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5102__A  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5096__B  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4945__B  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4758__A  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4623__D  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3648__A  (.DIODE(\MuI.a_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6174__A  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4783__B2  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4782__A  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4667__A1  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4666__B  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4468__A  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4467__B2  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4091__A  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3514__A  (.DIODE(\MuI.a_operand[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4667__B2  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4666__A  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4461__B  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4460__A1  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4208__B  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3492__A  (.DIODE(\MuI.a_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6148__A  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4343__B2  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4341__A  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4163__A  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4086__A  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3452__A  (.DIODE(\MuI.a_operand[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6151__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6041__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4298__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3957__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3868__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3791__A1  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3467__D  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3448__A  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3446__A  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3426__C  (.DIODE(\MuI.a_operand[25] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4728__A  (.DIODE(\MuI.a_operand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4424__A  (.DIODE(\MuI.a_operand[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5252__A1  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5196__B  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5113__B  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4956__A2  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4955__C  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4862__D  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4123__A  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3685__A  (.DIODE(\MuI.a_operand[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5000__D  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4826__D  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4782__D  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4666__D  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4461__D  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4460__B1  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4340__A  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4296__A  (.DIODE(\MuI.b_operand[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5231__B2  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5230__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4955__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4862__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4759__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4623__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3756__C  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3753__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3744__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3736__A  (.DIODE(\MuI.b_operand[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5844__A1_N  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5756__A  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5673__A  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4957__C  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4761__C  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4625__C  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3940__B  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3750__A  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3741__A  (.DIODE(\MuI.b_operand[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6116__B  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4972__C  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4711__C  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4515__A  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3883__A  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3696__A  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3657__A  (.DIODE(\MuI.b_operand[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3900__A  (.DIODE(\MuI.b_operand[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3540__A  (.DIODE(\MuI.b_operand[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5000__C  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4828__A2  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4826__C  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4782__C  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4666__C  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4461__C  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4460__A2  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4339__A  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4302__A  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4162__A  (.DIODE(\MuI.b_operand[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._6224__C  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4606__A  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4414__A  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4261__A  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3717__A  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3501__A  (.DIODE(\MuI.b_operand[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5152__B  (.DIODE(\MuI.b_operand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3866__A  (.DIODE(\MuI.b_operand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3795__A  (.DIODE(\MuI.b_operand[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._5250__A  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4947__D  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4848__D  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4750__D  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4643__B  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._4477__A  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_MuI._3771__A  (.DIODE(\MuI.b_operand[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A1 (.DIODE(\MuI.result[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(Operation[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(Operation[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(Operation[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(Operation[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__B2 (.DIODE(_00000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A2 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A2 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__D (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__A2 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__B (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__A2 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__C (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__B1 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__C (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__B (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__B (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__B (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A1 (.DIODE(_00011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__A (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B2 (.DIODE(_00012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__B2 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__B2 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__B2 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B2 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__A (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__A1 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__B (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__B (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A1 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__B1 (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__B (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__C (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__D (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B1 (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A2 (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__C (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__C (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__C (.DIODE(_00030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A2 (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__C (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A2 (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B1 (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A2_N (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__D (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__B1 (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__D (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__B (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B1 (.DIODE(_00033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B1 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A2 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__B1 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A2 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A2 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__D (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B1 (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__D (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__C (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A (.DIODE(_00035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__C (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A2 (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__D (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__B1 (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A2_N (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B2 (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A1 (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A2_N (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__D (.DIODE(_00036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__C (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__D (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__B1 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A2 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A2 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__D (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__B (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__B (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__B (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A1 (.DIODE(_00046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A2 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__C (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__B1 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B1 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__D (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A2 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__C (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B1 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A2 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__A2 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__C (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__B1 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__D (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A2 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__C (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B1 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B1 (.DIODE(_00048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B2 (.DIODE(_00049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__C (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__A (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A1 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A1 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__A (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A1_N (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A1 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A2 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__D (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__B (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A2 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A2 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B1 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A2 (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B (.DIODE(_00059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__B (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__B (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__B (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__B (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A1 (.DIODE(_00062_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__A (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__A (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B2 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__B2 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B2 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B2 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B2 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B1 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A2 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__B (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__B1 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A2 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A2 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__D (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__D (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A2 (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__D (.DIODE(_00072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__D (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__D (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__D (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A2 (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__D (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A2 (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__C (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A2 (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__A (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A2 (.DIODE(_00074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__C (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A1 (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__A (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A1_N (.DIODE(_00077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A1 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A1 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__B (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__B (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__A (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__A1 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__B (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A1 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__B (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A1 (.DIODE(_00081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__C (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__C (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__D (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A2 (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__C (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__D (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__C (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__D (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A (.DIODE(_00082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__D (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__D (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__B1 (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__C (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B1 (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__C (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__D (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B1 (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A2 (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A2 (.DIODE(_00083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__D (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__D (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__C (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__C (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__B1 (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__C (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__D (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A2 (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A (.DIODE(_00084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A2 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__C (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__D (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__D (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__B1 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A2 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B1 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A2 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B1 (.DIODE(_00085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__B2 (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B2 (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__B2 (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B2 (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A1 (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__C (.DIODE(_00088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__D (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__D (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__B1 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__B (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__B (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__B1 (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__C (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__C (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__D (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A (.DIODE(_00089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__C (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A2 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__B1 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__D (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__B1 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__B (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__D (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B1 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__D (.DIODE(_00090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A2 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__D (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__C (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__A2 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B1 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A2 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A1 (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__B (.DIODE(_00093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B2 (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A (.DIODE(_00095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__A1 (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A1 (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A1 (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B1 (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__B (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__B (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A2 (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B1 (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__D (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__D (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__C (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__B1 (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A2 (.DIODE(_00098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__C (.DIODE(_00105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(_00105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__C (.DIODE(_00105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__B2 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B2 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__B2 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A (.DIODE(_00124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__A (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__B (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__B (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__B (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__B (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A1 (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A1 (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A1 (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B (.DIODE(_00125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__B (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__B (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__B (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__B (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A1 (.DIODE(_00132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__A (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__A (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B2 (.DIODE(_00133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__C (.DIODE(_00141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B1 (.DIODE(_00141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__B (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__B (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__B (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__B (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__B (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__B (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__D (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12206__B (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__D (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B1 (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A2 (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A2 (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__C (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__B1 (.DIODE(_00153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__B (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A1 (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__D (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__B1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A2 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__B1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__B (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__B1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__C (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__D (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A2 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B2 (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__B (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__B1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__B (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__B (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B2 (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__A1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A1_N (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A1 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A1 (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A1 (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__A (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A1 (.DIODE(_00231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__B2 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__B2 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__B2 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B2 (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B1 (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__C (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__C (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A2 (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B1 (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A2_N (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__D (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__B1 (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__B (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A2 (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__D (.DIODE(_00259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A1 (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A1_N (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A1_N (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A1_N (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__C (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__C (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__B1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__C (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__A2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__B (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__D (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__D (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__C (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__D (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__D (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A2 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__C (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A1 (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A1 (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__C (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__C (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__B1 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__C (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__C (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__C (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__A2 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__C (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B1 (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__C (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__A (.DIODE(_00271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__C (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B1 (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A2_N (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__D (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__D (.DIODE(_00272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B2 (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__B2 (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__B2 (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B2 (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B2 (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(_00278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__B (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__B (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A1 (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__B (.DIODE(_00279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__B2 (.DIODE(_00281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A1 (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A1 (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A1 (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A1_N (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A1_N (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__C (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__C (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__D (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__C (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__D (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__D (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__C (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__D (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__A1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A1 (.DIODE(_00289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A1 (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__C (.DIODE(_00292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__B2 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__B2 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B2 (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__C (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A2 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__D (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A2 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__D (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A2 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A2_N (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B1 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__D (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__B (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B1 (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A2_N (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__D (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__D (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__D (.DIODE(_00303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__B (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A_N (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__A (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A1 (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A1 (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A1 (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A1 (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__A1 (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A (.DIODE(_00345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__C (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__B1 (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__C (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__B1 (.DIODE(_00363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__A2 (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__D (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__B1 (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__C (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__B1 (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A2 (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__D (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__B (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__C (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B (.DIODE(_00382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__B (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__C (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__D (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B1 (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__C (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__D (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A2 (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A2 (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B1 (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B1 (.DIODE(_00385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__D (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__B (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__C (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__B (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__C (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__C (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__D (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__B1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__C (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__C (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__D (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__B1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B2 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A1 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__D (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A2 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A2 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__B1 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__C (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A2 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__B (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__B (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B1 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__C (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__D (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__A2 (.DIODE(_00423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A1_N (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__A1 (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A1 (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__C (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A1 (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A1 (.DIODE(_00444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A1 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__C (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A2 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__D (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A2 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B1 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__C (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A2_N (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A2 (.DIODE(_00445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__B (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A1 (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A1 (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__B (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A1 (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__A (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__B (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A1 (.DIODE(_00462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B1 (.DIODE(_00471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07854__C (.DIODE(_00471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A (.DIODE(_00502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__A (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B2 (.DIODE(_00506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A2 (.DIODE(_00518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B (.DIODE(_00518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__B (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__B (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__B (.DIODE(_00519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__C (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__D (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__C (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B1 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__B (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A2 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__D (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A2 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__D (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B1 (.DIODE(_00530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__C (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A1 (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A2 (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__C (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__D (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__C (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__D (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__B1 (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A2_N (.DIODE(_00534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__B (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A1 (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__C (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__D (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__B (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A2 (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__B1 (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__D (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A2 (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A2_N (.DIODE(_00550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12194__B1 (.DIODE(_00555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__A1 (.DIODE(_00555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A1 (.DIODE(_00555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B2 (.DIODE(_00555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__B1 (.DIODE(_00555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12170__B1_N (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A1 (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A2 (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A2 (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B1 (.DIODE(_00566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A (.DIODE(_00567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__D (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A2 (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__D (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__C (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A2 (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__D (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__B1 (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__A2 (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__C (.DIODE(_00592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A1 (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B (.DIODE(_00596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A (.DIODE(_00610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A (.DIODE(_00610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B1 (.DIODE(_00617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__D (.DIODE(_00617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A2 (.DIODE(_00663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__C (.DIODE(_00663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A2 (.DIODE(_00663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A1 (.DIODE(_00664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__B (.DIODE(_00664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B1_N (.DIODE(_00664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__B_N (.DIODE(_00665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A_N (.DIODE(_00665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A1 (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A (.DIODE(_00672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__B (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__B (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11331__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__B (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A1 (.DIODE(_00676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__A1 (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A (.DIODE(_00691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__B1 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A1 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__B (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A1 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__C1 (.DIODE(_00702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A2 (.DIODE(_00702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A2 (.DIODE(_00702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__C (.DIODE(_00702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A (.DIODE(_00707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A (.DIODE(_00707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(_00707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__B (.DIODE(_00708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__B (.DIODE(_00708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B (.DIODE(_00708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__B (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A1 (.DIODE(_00727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B2 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A1 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A1 (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A (.DIODE(_00734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__B1_N (.DIODE(_00735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A2 (.DIODE(_00735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B (.DIODE(_00735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__B1 (.DIODE(_00739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__C (.DIODE(_00739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__D (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__D (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__B1 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__C (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__D (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A2 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B1 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__C (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__C (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__B1 (.DIODE(_00783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A2 (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__C (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A2 (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__D (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__C (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__D (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__A2 (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A2 (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__D (.DIODE(_00785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(_00810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A (.DIODE(_00810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__B (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__A (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B2 (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__B2 (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__B2 (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__B2 (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__A (.DIODE(_00877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__B (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A1 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__B (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08510__C (.DIODE(_00896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__B1 (.DIODE(_00896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__C (.DIODE(_00896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A1 (.DIODE(_00915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__A1 (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__B (.DIODE(_00919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A2 (.DIODE(_00919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__A (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__B2 (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__A (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__B2 (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__B2 (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__A (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B2 (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B2 (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__B (.DIODE(_00922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A2 (.DIODE(_00922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(_00923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B1_N (.DIODE(_00923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__B (.DIODE(_00929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B (.DIODE(_00929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A (.DIODE(_00934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A (.DIODE(_00934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(_00951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(_00951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__B (.DIODE(_00953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__B (.DIODE(_00953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B1 (.DIODE(_01026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__C (.DIODE(_01026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08465__A1 (.DIODE(_01071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A (.DIODE(_01071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(_01071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A (.DIODE(_01096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A (.DIODE(_01096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A_N (.DIODE(_01102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B (.DIODE(_01102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__B (.DIODE(_01140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__B (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__B (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__A (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__A (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B (.DIODE(_01150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__B (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A_N (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08554__B (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(_01203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A (.DIODE(_01203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__A (.DIODE(_01203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(_01203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__A (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__B (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__A1 (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__B (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__B (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A1 (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A1 (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A1 (.DIODE(_01206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__B1 (.DIODE(_01233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A (.DIODE(_01233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__C (.DIODE(_01266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B1 (.DIODE(_01266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__C (.DIODE(_01266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__B (.DIODE(_01325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__B (.DIODE(_01325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__B2 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__B2 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__B1 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A1 (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__B1 (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__B (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A2 (.DIODE(_01350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__B (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__B (.DIODE(_01378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__A (.DIODE(_01382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A (.DIODE(_01382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08774__B (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__B_N (.DIODE(_01387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08812__A (.DIODE(_01391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A (.DIODE(_01391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(_01394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__B (.DIODE(_01407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A1 (.DIODE(_01407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__A (.DIODE(_01407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A2 (.DIODE(_01409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08792__C (.DIODE(_01409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__A (.DIODE(_01419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A (.DIODE(_01419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08810__B (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__B_N (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A (.DIODE(_01427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__B (.DIODE(_01652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__C (.DIODE(_01668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__B1 (.DIODE(_01668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B1 (.DIODE(_01702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__A (.DIODE(_01702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__A1 (.DIODE(_01702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09167__A1 (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A (.DIODE(_01714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09165__B (.DIODE(_01722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B (.DIODE(_01722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__B (.DIODE(_01742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__B (.DIODE(_01742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__C1 (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B (.DIODE(_01881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__B1 (.DIODE(_01891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A1 (.DIODE(_01891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B1 (.DIODE(_01891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__B (.DIODE(_01891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__B (.DIODE(_01891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B1 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A2 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A2 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B2 (.DIODE(_01988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A (.DIODE(_02053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__A (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__B1 (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A (.DIODE(_02069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B2 (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B_N (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__A (.DIODE(_02096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__A (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B2 (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__A (.DIODE(_02107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__B2 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__B (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A1 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B2 (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__A (.DIODE(_02118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A1 (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A1 (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10069__B (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__A (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__A (.DIODE(_02129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__B (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A (.DIODE(_02194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__B (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__B2 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__B (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A (.DIODE(_02205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A1 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A1 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A1 (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__B (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A (.DIODE(_02216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__B (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__B (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__B (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__B (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A1 (.DIODE(_02229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__C (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A1 (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A (.DIODE(_02248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__B (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__B2 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A_N (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A1 (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A1_N (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__A (.DIODE(_02259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__A (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A1 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__B (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A_N (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__B_N (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__B2 (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__A1 (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A (.DIODE(_02334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B2 (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B2 (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A_N (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A1 (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__B1 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A1 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__B2 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_02350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__B (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A1_N (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A1 (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A1 (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A (.DIODE(_02377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B2 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__B_N (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A_N (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__B (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B2 (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__B2 (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B2 (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__B2 (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B2 (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__B2 (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B2 (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A (.DIODE(_02431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__B_N (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A_N (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__B2 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A1 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A1 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A1 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__A1 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__B (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A1 (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__A (.DIODE(_02474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__B (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__B (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A1 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A_N (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__B_N (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09432__B (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__A (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A1_N (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A1_N (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__C (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__A (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__A1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__A (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__B (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A_N (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A1 (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__A (.DIODE(_02550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__B2 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__B2 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__B2 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B2 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12510__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A1 (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A2 (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__A (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__B2 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A1 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A1 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A_N (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__B_N (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A1 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__B1 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__B2 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A1 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__B (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__B (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13390__A (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13296__A1 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__A1 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A1 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__A1 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__A2 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__A1 (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A1 (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A1 (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__B (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__A (.DIODE(_02647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__B (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__B (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A1 (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__A (.DIODE(_02658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A1 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A1 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__A (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__B (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__A (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__B_N (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__A1 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__A1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__A2 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__B (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13482__A (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__A1 (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__A (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13301__A1 (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__A1 (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__D (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__D (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__A (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A (.DIODE(_02705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13483__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__A1 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__B1 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__B1 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__B (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13451__C1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13243__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__A (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__B1 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A2 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__A (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__C (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__C (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__C (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__C (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__A (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13456__B1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__B1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__B1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__B1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__B1 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A3 (.DIODE(_02713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A2 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__A2 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A2 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A2 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B1 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A2 (.DIODE(_02719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B1 (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A (.DIODE(_02722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B2 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B_N (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A_N (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__A1 (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__A (.DIODE(_02723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A2 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__B1 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__B1 (.DIODE(_02724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13303__A2_N (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__B (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A2_N (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__B (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A2_N (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A2_N (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A2_N (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A2 (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__A (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__A (.DIODE(_02727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__B (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A2 (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A2_N (.DIODE(_02728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13397__A2 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A2 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B1 (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__A (.DIODE(_02731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__B1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__B1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__B1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A2 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B1 (.DIODE(_02732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__B1 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__B2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13300__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__B1 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__A2 (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A (.DIODE(_02738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__B1 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__A2 (.DIODE(_02739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13461__C1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13246__A (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__B (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__A (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__B1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__B1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A1 (.DIODE(_02741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__B1 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A2 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__B1 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A2 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A3 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A3 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A2 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A2 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A3 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A2 (.DIODE(_02745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13487__A1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13404__C1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__C1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__B1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A1 (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A (.DIODE(_02750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__B2 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13357__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13307__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A1 (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A (.DIODE(_02751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__A1 (.DIODE(_02752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__B2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__A (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__B_N (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__B2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__B2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__A (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__A (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__A (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A1 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__B2 (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__A (.DIODE(_02765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08742__A1 (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12887__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A2_N (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12879__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12878__A1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__C (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__A1 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__B2 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A1 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A1 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A_N (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__B_N (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A1 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__A1 (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__A (.DIODE(_02808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13427__A1 (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A1 (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__B2 (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13347__B (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__B1_N (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13312__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13311__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A1_N (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A1 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A1 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A1 (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A (.DIODE(_02840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12194__A1 (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B1 (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A1 (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__A (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B (.DIODE(_02848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A1_N (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A (.DIODE(_02851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A1 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__B2 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A2 (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A (.DIODE(_02860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__A (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A_N (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__B (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__A1 (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A (.DIODE(_02862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13406__A2 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A2 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13259__B (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__B (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A2 (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B2 (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__A (.DIODE(_02894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__B2 (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__B2 (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__A (.DIODE(_02905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__B2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__B_N (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__B (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A1 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__B2 (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A (.DIODE(_02916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13402__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13310__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13094__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__S (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12622__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__S (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__A2 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__B1 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11095__A2 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__B1 (.DIODE(_02931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__B2 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__B2 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11388__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__B2 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__A1 (.DIODE(_02935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13485__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A2 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11095__B1 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A2 (.DIODE(_02938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__A2 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A2 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A2 (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A2_N (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__B (.DIODE(_02941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13299__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B1 (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A (.DIODE(_02944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A2 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__B1 (.DIODE(_02945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__B (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A1 (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06770__A (.DIODE(_02948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__B (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__B (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__B (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__B (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__B (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A1 (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__A (.DIODE(_02959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A1 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A1 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A1 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B2 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A_N (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A1 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__A (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A1 (.DIODE(_02977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__A (.DIODE(_02977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__B (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__B (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__A1 (.DIODE(_02980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__B2 (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B2 (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__B2 (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__B2 (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A (.DIODE(_02983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A1 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A1 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A1 (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__B (.DIODE(_02984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A1 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__B1 (.DIODE(_02991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A (.DIODE(_02999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__B (.DIODE(_02999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A1 (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__A1 (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__A (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08637__C (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1_N (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__C (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A1_N (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A (.DIODE(_03002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__A1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A1 (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A1 (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__A_N (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__B_N (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A1 (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A1 (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A1 (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A (.DIODE(_03024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A2 (.DIODE(_03046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A (.DIODE(_03046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A2 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__B1 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__C (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A2 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__B (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B1 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__B (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__B (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A2 (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__D (.DIODE(_03047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A2 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A2 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A2 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__B1 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__C (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A2 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__B (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__C (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__D (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__B1 (.DIODE(_03051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__B (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A_N (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__B2 (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__B2 (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A (.DIODE(_03067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__B1 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12743__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__B (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__B1 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__B (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__D (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__D (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__B (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A2 (.DIODE(_03071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__B (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A1 (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A (.DIODE(_03099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A1 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__B2 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A_N (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A1 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__B (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__A1 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__B (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A_N (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__B (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__B1 (.DIODE(_03119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13419__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13233__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__B1 (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A (.DIODE(_03133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__C1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13306__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__B1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__B1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A1 (.DIODE(_03134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A (.DIODE(_03152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__A1 (.DIODE(_03157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A (.DIODE(_03157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A1 (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__C (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__C (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__C (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A (.DIODE(_03163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__B2 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A1 (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A1_N (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__C (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A1_N (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__A (.DIODE(_03174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__A2 (.DIODE(_03186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__A_N (.DIODE(_03186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__B1_N (.DIODE(_03186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__A (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__B2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__B2 (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__A (.DIODE(_03228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__B2 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A1 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__B_N (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A_N (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__B2 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B2 (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__A (.DIODE(_03239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__C (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__B1 (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A2 (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__B (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__D (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A2 (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__B (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__B (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__C (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__D (.DIODE(_03247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__B1 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12628__B (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A2 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__B (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B1 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A2 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__B (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__B (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__A2 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__B (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__B (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A1 (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A (.DIODE(_03271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A1 (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__A (.DIODE(_03282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A2 (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__B (.DIODE(_03289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__B_N (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__B2 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A_N (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__B (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A1 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__C1 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__B2 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__B2 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A1_N (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__B1 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__B2 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A1_N (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A1_N (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__B (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__B2 (.DIODE(_03306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__A1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__B1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12873__B1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__C1 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A2 (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__A (.DIODE(_03314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A1 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A1 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__B2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__B1 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__A1 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11097__A2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__A2 (.DIODE(_03315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A1 (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__A (.DIODE(_03324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__B1 (.DIODE(_03330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__A (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A (.DIODE(_03331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A1 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A1 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A1_N (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A1_N (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__A (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__B2 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A1_N (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B_N (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A_N (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A1 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12741__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B2 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__A (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__B2 (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B2 (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B2 (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A (.DIODE(_03389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__A (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A1 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A1 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A1 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__B (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A_N (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A1 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B1 (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A (.DIODE(_03400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__C (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12661__A2 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__D (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__B1 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A2 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__A2 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__C (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__D (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__B (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A2 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__C (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A2 (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__A2 (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__C (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__D (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B1 (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__C (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__D (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B1 (.DIODE(_03425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__B (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A1 (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__A (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A1 (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A1 (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__B (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__B (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__B (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A1 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__A (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12630__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__C (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__B (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__B1 (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A2 (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__C (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__B1 (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A2 (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__C (.DIODE(_03444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__B1 (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__D (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__C (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__B1 (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__B (.DIODE(_03449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__B2 (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__A (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__B2 (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A1 (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__B (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A_N (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B_N (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A1 (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__B (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A (.DIODE(_03454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__B (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__B (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13295__C1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__A1 (.DIODE(_03489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__B1 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A1 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__A (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__B1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__B_N (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A_N (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__A (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A (.DIODE(_03509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__A1 (.DIODE(_03509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A (.DIODE(_03534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__A (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__B2 (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__A (.DIODE(_03550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A1 (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A1 (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__B2 (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B2 (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A1 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__B (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A1 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__B (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__A1 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A1 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A1 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__B (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__B_N (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__B2 (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__B (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A1 (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__A (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__A (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A_N (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A (.DIODE(_03626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__B (.DIODE(_03655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__B (.DIODE(_03655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__A1 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A1 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__A (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A1 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__A1 (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__A (.DIODE(_03669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__B1 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A2 (.DIODE(_03675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__B2 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13317__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__A1 (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__B_N (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__A_N (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__B (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__A (.DIODE(_03680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A1 (.DIODE(_03692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__B1 (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__A (.DIODE(_03713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__C (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B1 (.DIODE(_03717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A (.DIODE(_03722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A1 (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__A (.DIODE(_03733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A1 (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A1 (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__A1 (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__A (.DIODE(_03744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A1 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__A1 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__A1 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__A (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A3 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B1 (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__C (.DIODE(_03762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__A (.DIODE(_03798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A1 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A1 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A1 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__A1 (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__A (.DIODE(_03809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A (.DIODE(_03820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__A2 (.DIODE(_03828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__B (.DIODE(_03828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__A (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__A (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A1 (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A (.DIODE(_03831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A1 (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__A (.DIODE(_03842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A2 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__B (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__C (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A2_N (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__D (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A2_N (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__D (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__C (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A2 (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__A (.DIODE(_03873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__B1 (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__A (.DIODE(_03879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A2 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__C1 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__B (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__C (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__D (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__C (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08547__A2 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__B (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A2 (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__A (.DIODE(_03884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__B (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__B (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A2 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__A2 (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A2_N (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__C (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__C (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A (.DIODE(_03895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__A_N (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__A2 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A2 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A2 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08551__A2 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__C1 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A2 (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A (.DIODE(_03906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A1_N (.DIODE(_03913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A (.DIODE(_03913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__C (.DIODE(_03913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B_N (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A2 (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__B (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A2 (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__C1 (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09684__A2 (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__B (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__B (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__A (.DIODE(_03917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__B2 (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A2 (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A1_N (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A2 (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__B (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__B (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__A (.DIODE(_03928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__A (.DIODE(_03939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__D (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__B (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B1 (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A2 (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A2 (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__C (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__C (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A2 (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__B1 (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A2 (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__D (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__B (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__D (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A2 (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__B (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__D (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A2_N (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__B (.DIODE(_03973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__B1 (.DIODE(_03973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B1 (.DIODE(_03973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__A (.DIODE(_03974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A2 (.DIODE(_03974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B2 (.DIODE(_03974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__B (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09879__A2_N (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__B1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__B1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A2 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__D (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A2 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B1 (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__A (.DIODE(_03982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A_N (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B_N (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09646__B1 (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09187__A2 (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__B1 (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__D (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__D (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__A (.DIODE(_03993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A2 (.DIODE(_04000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__B (.DIODE(_04000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B1 (.DIODE(_04002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B2 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A2 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A2 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__A (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__B1 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A2 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A1 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B1 (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__A (.DIODE(_04004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__C1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__B2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__B2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B2 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__B1 (.DIODE(_04011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A (.DIODE(_04015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A2 (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A2 (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A2_N (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__D (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__D (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B1 (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__C (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A2 (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__D (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__B (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__B1 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__C (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A2_N (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A2_N (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__A (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__B (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A2 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A2 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A2 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A2 (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A2_N (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__B (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A (.DIODE(_04057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__B2 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A_N (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A2 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A1 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A2 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__B (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__B (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B2 (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__A (.DIODE(_04068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__B1 (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A1 (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__B (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11312__A2 (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__B (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__D (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A2 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A2_N (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__D (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__D (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__C (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A2 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__B (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__B1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__A (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B1 (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A_N (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__B (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A2_N (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A2 (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B1 (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A2_N (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A2 (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__B2 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A2 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A2 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A1 (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__B (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__B (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__A (.DIODE(_04133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__A (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A2 (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B (.DIODE(_04149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__B1_N (.DIODE(_04151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__B1 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__A1 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A2 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__A2 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B1 (.DIODE(_04159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13400__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__B1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A1 (.DIODE(_04161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__B (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__B (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__D (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__D (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A2 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__C (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__A (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__D (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A2 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__A (.DIODE(_04176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__B (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A_N (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A2 (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__B (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A2_N (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A (.DIODE(_04186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__B2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B_N (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A1_N (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A2 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A1 (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__B (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__B (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__B (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A (.DIODE(_04197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A (.DIODE(_04208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A1 (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12955__B1 (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__B1 (.DIODE(_04211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__B (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__D (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__D (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__B (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__D (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__B1 (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__D (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__D (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__B1 (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__B1_N (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B (.DIODE(_04233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__B1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__C (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A2 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__C (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__C (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A2 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__D (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__B (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__B (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__B (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A_N (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A2 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A2_N (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A2 (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A2_N (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A (.DIODE(_04251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__B2 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__B (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A1_N (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__B (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__B (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__A (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__B1 (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(_04269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A (.DIODE(_04273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B1 (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A2 (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__C (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__C (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__B (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A2 (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__D (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__C (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__A (.DIODE(_04302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__A1 (.DIODE(_04302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__B (.DIODE(_04302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__A2 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__C (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__D (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A2 (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__B (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A2_N (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__B1 (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__D (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__D (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B1 (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__B1 (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A (.DIODE(_04305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__B1 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__B (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A2 (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__B (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A2 (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A2_N (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A2_N (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A2 (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__B (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__A (.DIODE(_04316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__A (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B2 (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A1_N (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A2 (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__A2 (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__B2 (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A (.DIODE(_04338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__C (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__C (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__C (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A2 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A2 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__C (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B1 (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__B1 (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A2 (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__D (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B1 (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A2_N (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__D (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A2 (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A2_N (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__B (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A1 (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A (.DIODE(_04369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__B (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A2 (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__B (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__A2 (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A2_N (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__B2 (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__A (.DIODE(_04380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__B2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__B (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A1_N (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B2 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__B (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__B_N (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__A (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A (.DIODE(_04413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__B1 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A2 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A2 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__B (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B1 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A2 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__D (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__C (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__A (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__C (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__B (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__B (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A2 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__B (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__B1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__C (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__A (.DIODE(_04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__B1 (.DIODE(_04446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A (.DIODE(_04446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__B (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__A2 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__B (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__B1 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__B (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A2 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A2 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B2 (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__A (.DIODE(_04456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__B2 (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A2 (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1_N (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__B (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A1 (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__B (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A_N (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A (.DIODE(_04467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__A (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__A1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__B1 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__A2 (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__C1 (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__A (.DIODE(_04489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__C1 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__B1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A2 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A2 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__C (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A2 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__C (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__C (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__D (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__B1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__C (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A2 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__D (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__B1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A2_N (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A2_N (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__D (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__B (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__A2 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__B (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__B (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A2 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08727__A2 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A2 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__B (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__B2 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A2 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A1_N (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__B2 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__B1 (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__A (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__D (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__B (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__D (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__D (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__C (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__B1 (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__B (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A2 (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A (.DIODE(_04574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__B (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__D (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A2 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__C (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__B (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__C (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B1 (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A (.DIODE(_04585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A2 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__B2 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A1 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A2 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A2 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A1 (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__B1 (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__A (.DIODE(_04604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__A (.DIODE(_04606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A (.DIODE(_04606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__B2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__A1_N (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B2 (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__B_N (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B1 (.DIODE(_04623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__B1 (.DIODE(_04631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12888__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12524__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__S (.DIODE(_04635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B1 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A2 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__B1 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A2 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A2 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__D (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__D (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A2 (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A (.DIODE(_04638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A2 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A2 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__B1 (.DIODE(_04642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__C (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A2 (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__B1 (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__C (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__B (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__B (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__B1 (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__C (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__D (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__A (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__B (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A2 (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__B (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__B2 (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A2 (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A2 (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A2 (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__A (.DIODE(_04660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__B2 (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__B (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A2 (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A1 (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__B2 (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A_N (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__A (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A (.DIODE(_04671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__A2 (.DIODE(_04677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A (.DIODE(_04677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__A1 (.DIODE(_04677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__A1 (.DIODE(_04678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A (.DIODE(_04678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__A2 (.DIODE(_04678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__B1_N (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__A2 (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__B (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__B (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__D (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__D (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__C (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A2 (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B1 (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__C (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__D (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A (.DIODE(_04703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__D (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__B (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__C (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A2 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__D (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B1 (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A2_N (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__B (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__D (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__B1 (.DIODE(_04721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__A (.DIODE(_04721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__B (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__B (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A2 (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__B (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B2 (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A1 (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__B (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A2 (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__A2_N (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A (.DIODE(_04725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__B2 (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A1_N (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A2 (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11907__B (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A1 (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__B_N (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__B (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A (.DIODE(_04736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A1 (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__B1 (.DIODE(_04755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A2 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__C1 (.DIODE(_04756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__B (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A2 (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__C (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__B (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__C (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A2 (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__B1 (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A2 (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__D (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__A (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__C (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__D (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__B (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A2 (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__D (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__B (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__B (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B1 (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__D (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__A (.DIODE(_04789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__A1_N (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__B2 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__B (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__B (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__B2 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__B (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A1 (.DIODE(_04803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__A (.DIODE(_04803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__B1 (.DIODE(_04803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__B1 (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__B1 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A2 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__B1 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A2 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A2 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__D (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B1 (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__C (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A (.DIODE(_04832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__B1 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__D (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__B (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__A2 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B1 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__D (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__C (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A2 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__B (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__B (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A2 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__B (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__B2 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__B (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A2 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A2 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__B1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A1 (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__A (.DIODE(_04864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__B2 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__B (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A1_N (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__A2 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A2 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__B2 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__B (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A_N (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__A (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A2 (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__B (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__B1 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B1 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B1 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B1 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A2 (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__C (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__C (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__D (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A (.DIODE(_04896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A2 (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B1 (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__C (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A2 (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__B1 (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__B (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__D (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B1 (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__D (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A (.DIODE(_04907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__A2 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__B2 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A2 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A2 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B2 (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A2 (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A1_N (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B2 (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A_N (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__B_N (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(_04929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__B1 (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A2 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__C (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A2 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__B1 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__B1 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__D (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A2 (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(_04961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__C (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A2 (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__D (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__B1 (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__C (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__D (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__B1 (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__B (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A2_N (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(_04972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__B (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12367__A2 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__B (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A2 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__B2 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__B (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__A2 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__B (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A1 (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A (.DIODE(_04983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A1 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__B1 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__A2 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__C1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__B (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B2 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A2 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__A2 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12504__A1_N (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A2 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A1 (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__A_N (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__A2 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__C (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__C (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A2 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__B1 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A2 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__B (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__C (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A2 (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(_05025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__C (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A2 (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__B1 (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__C (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__D (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A2 (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A2_N (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__D (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B1 (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A (.DIODE(_05036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A (.DIODE(_05041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__C (.DIODE(_05041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A2 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__B2 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A2 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__A2 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__A2 (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12220__A (.DIODE(_05052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__B2 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__B (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A2 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__B2 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__B (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10170__A (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__A (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A1 (.DIODE(_05092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__B1 (.DIODE(_05092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__A (.DIODE(_05092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__A2 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__B1 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__D (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A2 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__D (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__C (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__D (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A (.DIODE(_05101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A2 (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__B1 (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B1 (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__C (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__A (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B1 (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B1 (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__D (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_05112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12575__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__B2 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__A2 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__B2 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A1 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__A (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__B1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__B1 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A2 (.DIODE(_05127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__C1 (.DIODE(_05127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__B2 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A_N (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__B (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A1 (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__B (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__B (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__B (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A (.DIODE(_05134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__B1 (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__B (.DIODE(_05160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B1 (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__C (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A2 (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__D (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__C (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__D (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__C (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__C (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__B (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__C (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__A2 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__C (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A2 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__D (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__B1 (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__A (.DIODE(_05187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12568__A2 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__B (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__B (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__B1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__D (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__B1 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__B (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A2 (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A (.DIODE(_05198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__B2 (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__B (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1_N (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__B2 (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__B (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__B (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__B (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A_N (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(_05209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__B1_N (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__C_N (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A1 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A2 (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__B (.DIODE(_05233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__C (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__B1 (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__C (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A2 (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__D (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__C (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__D (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__B1 (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__C (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A2 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__D (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__C (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__D (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__D (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__B1 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__C (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A2 (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A (.DIODE(_05252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__B (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__B (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__A2 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12566__B (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__B (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A2 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__B (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A2 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A2 (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(_05262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__B1 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12489__A1 (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__A2 (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__B2 (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A2 (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A1_N (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__A2 (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__B2 (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__B (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A (.DIODE(_05273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__D (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__D (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A2 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__C (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B1 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__B1 (.DIODE(_05308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A (.DIODE(_05308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__D (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__D (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A2 (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__A2 (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__C (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__B1 (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__B (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(_05316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__B (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A2 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__B1 (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A (.DIODE(_05327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__B (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B2 (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A1 (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12941__A2 (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12881__A1 (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__A (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__B (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A (.DIODE(_05338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__B1 (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A1 (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A1 (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A2 (.DIODE(_05341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__B (.DIODE(_05341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B1 (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__C (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A2 (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__D (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__D (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A2 (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__C (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A (.DIODE(_05370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12518__B1 (.DIODE(_05376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__C1 (.DIODE(_05377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A2 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A2 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__B (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B1 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__B1 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__C (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A2 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__D (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B1 (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A (.DIODE(_05380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A2 (.DIODE(_05387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12927__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12581__A2 (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__C (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A2 (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A (.DIODE(_05391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B2 (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__A (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A2 (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__A1_N (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A2 (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__A1 (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__A_N (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__B (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__A (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A (.DIODE(_05402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B1 (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__D (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__C (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A2 (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__C (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A2 (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__D (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A2 (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A2 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__B1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__C (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__B1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__B1 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__C (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__D (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__A2 (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__B (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__A (.DIODE(_05445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12923__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12216__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__B (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__A2 (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(_05456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A1 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__B (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A1 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13084__A2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__B2 (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__B (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A (.DIODE(_05467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__A (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__B1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12612__A2 (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__C1 (.DIODE(_05476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__D (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A2 (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__D (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__D (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A2 (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A2 (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__C (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A (.DIODE(_05498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__C (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__B1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__C (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__C (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__D (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__D (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A2 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__B1 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A2 (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A (.DIODE(_05509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A2 (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A2 (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__B (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__A2 (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__A (.DIODE(_05520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13241__B (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13236__B2 (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A2 (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A2 (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A1_N (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A1 (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__A_N (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__B (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A (.DIODE(_05531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12787__A1 (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__B1 (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A1 (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__B1 (.DIODE(_05559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__C (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A2 (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__B1 (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__C (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__D (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B1 (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A2 (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B1 (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A (.DIODE(_05563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__D (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__D (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__C (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B1 (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B1 (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__C (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__B1 (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_05574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__B1 (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A2 (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13058__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__C (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__A2 (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__B (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A (.DIODE(_05585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13299__B2 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13237__B (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13235__A1 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B2 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A2 (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__B (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__B (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__D (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__D (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__A (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__C (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__D (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__D (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__B1 (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A2 (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__B1 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10874__C (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A2 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A2 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__B1 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__D (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A2 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__B1 (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A (.DIODE(_05638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12917__D (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__C (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A2 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A2 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13215__A2 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__B (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__A2 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__B (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__C (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12916__B1 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__B (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__A2 (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(_05660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__B2 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13303__A1_N (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13239__A1 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__B (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__B (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__B (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__B (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__B1 (.DIODE(_05676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A1 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__A (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__B1 (.DIODE(_05700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__A2 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A2 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__C (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__B1 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A2 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__D (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__A2 (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__D (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__B (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A (.DIODE(_05702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13273__B (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13210__A2 (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__B (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__A2 (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__B (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A2 (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__D (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A2 (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__B (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A (.DIODE(_05713_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__B2 (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13351__A2 (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A1_N (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13337__A2 (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13302__A1 (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A2 (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__B (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__B (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A (.DIODE(_05724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__B1 (.DIODE(_05754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__D (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__C (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A2 (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__C (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__B1 (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__B (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__C (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A2 (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B1 (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A (.DIODE(_05756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12953__C (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12952__A2 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__A1 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12885__A2 (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A2 (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__B1 (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__D (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A2_N (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__C (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__D (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B1 (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A2 (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11454__B1 (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__A (.DIODE(_05767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13268__A2 (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__B (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13115__B (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__B1 (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A2 (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__A2 (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__B (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__B (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__A (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__A (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13353__B2 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13329__B (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13267__B (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__B (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__B (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__B1 (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A2 (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__B1 (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__D (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A2 (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__C (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__B1 (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__D (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__A (.DIODE(_05820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A2 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__D (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A2 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A2 (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__B (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A2 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__B (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13261__B (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A2 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13133__A2 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__B (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__A2 (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A2_N (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(_05842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B1 (.DIODE(_05845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__B2 (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13433__A (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A1 (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13412__A2 (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13394__B2 (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__B (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A_N (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__A (.DIODE(_05853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__B (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13388__A1 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13120__B (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__A2 (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__B1_N (.DIODE(_05883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__B1 (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__B (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__C (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__B1 (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__D (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B1 (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__B (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__D (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__B (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A (.DIODE(_05884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__B1 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A2 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A2 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__C (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__B2 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A1 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A2 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__B (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A2 (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A (.DIODE(_05895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A2 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__C (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__B1 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__B (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__A2 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A2 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__A2 (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__B (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__B (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A (.DIODE(_05906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13484__B2 (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13465__A (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A2 (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__B2 (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__B (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(_05917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A2 (.DIODE(_05925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__C (.DIODE(_05925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__B1 (.DIODE(_05925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__B2 (.DIODE(_05926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__D (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__B1 (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__B1 (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__D (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A1 (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A (.DIODE(_05948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A2 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__B1 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B1 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__B (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__B (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__B2 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B1 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__B (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__B2 (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__B (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__B (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__B (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__D (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__A1 (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__B (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A2 (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__B (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B1 (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__A (.DIODE(_05970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__B1 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13317__B (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13316__D (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A2 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13134__B1 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A2 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__B1 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__B (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11952__B1 (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(_05981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13481__A1_N (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13464__A1 (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13407__B (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__B (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A2 (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__C1 (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__B (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__B (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(_05992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__B1 (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__B (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A2 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A3 (.DIODE(_06000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__A (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__B2 (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__B (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__A (.DIODE(_06016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A2 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13238__A2 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A2 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A2 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__B1 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__B1 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__B1 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13398__A2 (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12884__A2 (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A2 (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A2 (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__B1 (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A (.DIODE(_06056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__C (.DIODE(_06091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13247__B1 (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13249__A (.DIODE(_06157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A2 (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13305__A3 (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13355__A2 (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__B (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A2 (.DIODE(_06305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13399__A3 (.DIODE(_06306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A2 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__A (.DIODE(_06376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A2 (.DIODE(_06394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A3 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13494__A (.DIODE(_06408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__B1 (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__B (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__A (.DIODE(_06427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13469__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13387__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__B1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__A (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__A1 (.DIODE(_06428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11337__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(_06429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A2 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__D (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__C (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__D (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__C (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A2 (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__C (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__D (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__D (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__C (.DIODE(_06430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__D (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__D (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__B1 (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__D (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__C (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__C (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__C (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__D (.DIODE(_06431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B1 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__B (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__C (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__A (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__D (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__B1 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__D (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__D (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__A2 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A2 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__C (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__D (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__C (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__C (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A2 (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__A (.DIODE(_06436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__B (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__C (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__B1 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A2_N (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08802__B (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__A2 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A2 (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__D (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A2_N (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__D (.DIODE(_06437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A1_N (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__C (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A1_N (.DIODE(_06439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__B (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__B (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__B (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(_06442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__B (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__B (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A2 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__B1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__B (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__D (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__D (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__D (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B1 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B2 (.DIODE(_06444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__B (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09640__B1 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__B1 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__D (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B1 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__C (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__D (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A2 (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__D (.DIODE(_06446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(_06452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A (.DIODE(_06455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__B (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09199__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__C (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__D (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__A (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A2 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__C (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__D (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__D (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__B1 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A2 (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B (.DIODE(_06461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__B (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A1 (.DIODE(_06463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__C (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__D (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__D (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A2 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__B1 (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__D (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__B (.DIODE(_06466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__B2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09314__B2 (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_06469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__A1 (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B1_N (.DIODE(_06470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__C (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__C (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__D (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__C (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__C (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__B (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__C (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__D (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A2 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__B1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__B (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A2 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12257__D (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__B1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__B1 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__B (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A2 (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__B (.DIODE(_06477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__B2 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__B2 (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A (.DIODE(_06479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__A1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A1 (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B (.DIODE(_06480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__A (.DIODE(_06488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__C (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__C (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11616__D (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__C (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__D (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B1 (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__B (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A1 (.DIODE(_06491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__A (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__B2 (.DIODE(_06492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__B2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A1 (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B (.DIODE(_06495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__B (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__B (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A1 (.DIODE(_06500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B2 (.DIODE(_06501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__B2 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__B2 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B2 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B2 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__A (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__B (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__B (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A1 (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__B (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__B (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__B (.DIODE(_06504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A1 (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__B (.DIODE(_06513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__B (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__B (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A1 (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__B (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A (.DIODE(_06515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__B (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__B (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__B (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A1 (.DIODE(_06516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__D (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__B (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__D (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__C (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__B1 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__A2 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A2 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B1 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A2 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__D (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__C (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B1 (.DIODE(_06518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__B2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B2 (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A (.DIODE(_06519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__C (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__D (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__B1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__C (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__D (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__A2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__B (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__B (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__B (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B2 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__C (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__C (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__D (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__C (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A2 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10874__D (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A2 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__B1 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A2 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A1_N (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__C (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09424__C (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__A (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A1_N (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A1_N (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A1 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__D (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B1 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__B1 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__C (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A2 (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A1 (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A1 (.DIODE(_06558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A (.DIODE(_06558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A1 (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A1 (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A1 (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A2 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A2 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__B1 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__B (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A2 (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__B (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__C (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__B (.DIODE(_06561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__C (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A2 (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11308__B1 (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__A2 (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__D (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__B (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__C (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__D (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__C (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A2 (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09434__B2 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__B2 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__B2 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__B2 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B2 (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A (.DIODE(_06564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B2 (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A (.DIODE(_06565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A2 (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__D (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11434__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__D (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B1 (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B1 (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__D (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__B1 (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A2 (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B2 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B2 (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08896__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(_06578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__A1 (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__B (.DIODE(_06579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__B (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__C (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A2 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__C (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__D (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B1 (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__D (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__C (.DIODE(_06580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__D (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__D (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__B1 (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A2 (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08604__C (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B1 (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__C (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__D (.DIODE(_06581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10874__B (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__B (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__B (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A1 (.DIODE(_06583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__B1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__D (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__B1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__A2 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__D (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A2 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__C (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B1 (.DIODE(_06584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10874__A (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B2 (.DIODE(_06585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__B1 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__D (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__C (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__C (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A2 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__D (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B1 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A2 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B1 (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__D (.DIODE(_06591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__A (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A1_N (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A1_N (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__A1_N (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__C (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A1_N (.DIODE(_06593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B2 (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__A (.DIODE(_06598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10701__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A1 (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(_06599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__B (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__B (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A1 (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__A1 (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A1 (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__B (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A1 (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__B (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A1 (.DIODE(_06601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__B1 (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A2 (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__C (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__D (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__C (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__B (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__C (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__D (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__D (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A (.DIODE(_06602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A2 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__C (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__B1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__C (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__B (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__D (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B1 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A2 (.DIODE(_06603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__B1 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A2 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__D (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__B (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__C (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__D (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__B (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A2 (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__D (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A (.DIODE(_06604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A2 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__C (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__C (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10844__D (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__B (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__C (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A2 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B1 (.DIODE(_06605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__B2 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08467__B2 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B2 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B2 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B2 (.DIODE(_06606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__C (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__C (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__C (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__C (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__A (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__C (.DIODE(_06608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A1 (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__A1 (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A1_N (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A1_N (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__A1_N (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A1 (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A1_N (.DIODE(_06610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__B1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A2 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__C (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B1 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__D (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__C (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A2 (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__C (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A (.DIODE(_06611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A2 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__C (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__B1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A2 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__B1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__C (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A2 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__B (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B1 (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A (.DIODE(_06612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A2 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__B (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A1 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__B (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__A2 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__B1 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A2 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__B (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A2_N (.DIODE(_06613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__A1 (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A1_N (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__C (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A1_N (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A1_N (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A1 (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A1_N (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A1_N (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__B (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08897__A1 (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A1 (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A1 (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A1 (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A1 (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__B (.DIODE(_06622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__B1 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__B (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__C (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__D (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B1 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__B1 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A2 (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__C (.DIODE(_06623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B1_N (.DIODE(_06629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A1 (.DIODE(_06629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A (.DIODE(_06629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__B (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__B (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A1 (.DIODE(_06630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__A (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B2 (.DIODE(_06631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B (.DIODE(_06635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B (.DIODE(_06635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A1_N (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__C (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__C (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A (.DIODE(_06663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__C (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__D (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A2 (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__D (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__B (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A2 (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__A2 (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B1 (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__B (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__D (.DIODE(_06666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A1_N (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A1_N (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__C (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__C (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__C (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A (.DIODE(_06680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__B2 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__B (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09454__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__B (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A1 (.DIODE(_06682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(a_operand[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(a_operand[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(a_operand[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(a_operand[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(a_operand[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(a_operand[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(a_operand[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(a_operand[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(a_operand[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(a_operand[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(a_operand[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(a_operand[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(a_operand[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(a_operand[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(a_operand[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(a_operand[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(a_operand[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(a_operand[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(a_operand[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(a_operand[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(a_operand[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(a_operand[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(a_operand[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(a_operand[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(a_operand[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(a_operand[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(a_operand[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(a_operand[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(a_operand[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(a_operand[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(a_operand[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(a_operand[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(b_operand[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(b_operand[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(b_operand[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(b_operand[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(b_operand[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(b_operand[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(b_operand[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(b_operand[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(b_operand[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(b_operand[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(b_operand[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(b_operand[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(b_operand[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(b_operand[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(b_operand[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(b_operand[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(b_operand[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(b_operand[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(b_operand[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(b_operand[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(b_operand[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(b_operand[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(b_operand[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(b_operand[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(b_operand[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(b_operand[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(b_operand[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(b_operand[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(b_operand[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(b_operand[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(b_operand[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(b_operand[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06693__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__B_N (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06683__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1030__A3  (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0928__A0  (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__C (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1252__A0  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1014__A1  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0867__A2  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0863__A2  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0859__B2  (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__D (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1266__A0  (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1012__A1  (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0854__A  (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1277__A0  (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1004__A1  (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0850__A  (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1294__A0  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1002__A1  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0853__B2  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0852__B2  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__C (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__D (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1308__A0  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1008__A1  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0853__A2  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0849__B2  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__D (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1322__A0  (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1006__A1  (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0855__A_N  (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0849__A2  (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1331__A0  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0960__A1  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__D (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1347__A0  (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0958__A1  (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0825__A2  (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0817__B  (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__C (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__C (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1356__A0  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0969__A1  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0822__B  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0820__B2  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1367__A0  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0967__A1  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0821__B  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0820__A2  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1088__A0  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1071__A3  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1030__A1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__C (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1374__A0  (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0974__A1  (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0807__A  (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__D (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1386__A0  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0972__A1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0806__A  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1396__A0  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0989__A1  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0814__C_N  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0812__B  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__C (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0930__A  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0907__A0  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0805__A  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0933__A  (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0884__A  (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0881__A  (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0936__A1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0915__A0  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0879__A  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0878__B_N  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__C (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0943__A1  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0917__A0  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0888__B1  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0877__B  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0948__A1  (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0954__A1  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0923__A0  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1113__A0  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1071__A1  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1031__A3  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0837__A  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__C (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__D (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0910__B_N  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0900__B  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0896__A  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0895__A  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__D (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1675__A1  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1043__A  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0927__A  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1137__A0  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1073__A3  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1031__A1  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1153__A0  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1073__A2  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1171__A0  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1189__A0  (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1025__A1  (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__C (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07471__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1210__A0  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1026__A1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0861__A2_N  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0835__A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1224__A0  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1016__A1  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0860__A  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1241__A0  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1017__A1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0867__B2  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0864__B2  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0863__B2  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1030__A2  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0928__A1  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0839__B  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1252__A1  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1014__A0  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0858__A  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1277__A1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1004__A0  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0856__A2  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0852__A2_N  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1294__A1  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1002__A0  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0851__A  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1308__A1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1331__A1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0960__A0  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0824__A  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1356__A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1367__A1  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0967__A0  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1088__A1  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1071__A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1374__A1  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0974__A0  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0874__A1  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0808__B1  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1386__A1  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0972__A0  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0813__A1  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0808__A1  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1396__A1  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0989__A0  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0814__A  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0812__A  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0929__B1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0932__B1  (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0936__A0  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0915__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0879__B_N  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0878__A  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0943__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0917__A1  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0889__A2_N  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0877__A  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0946__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0919__A1  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0887__A  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0948__A0  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0921__A1  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0894__A1  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0890__A  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__C (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0954__A0  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0923__A1  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0898__B_N  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0893__A  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1113__A1  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1071__A0  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1031__A2  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0910__A  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0900__A_N  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0896__B  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0895__B  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0926__B  (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1137__A1  (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1073__A1  (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1153__A1  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1073__A0  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1171__A1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1067__A0  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1189__A1  (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1210__A1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1026__A0  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0833__A  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1224__A1  (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1016__A0  (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1241__A1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1017__A0  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0862__A  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0864__A2_N  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0861__B2  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1025__A0  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0834__A  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0827__B  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1028__A0  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0830__A  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0828__B  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1028__A2  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0844__B  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0831__A  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1031__A0  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0845__A1  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0843__A1  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0843__B1  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0841__A1  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0876__A  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0911__A  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0885__A2  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0881__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0907__A1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0815__A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0810__B  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0809__B  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__C (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0839__A_N  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A2_N (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__C (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1030__A0  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0840__B  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0838__A  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0818__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0969__A0  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0819__A  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1347__A1  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0958__A0  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0816__A  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1322__A1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1006__A0  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0855__B  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0847__A  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1008__A0  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0848__A  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__C (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1266__A1  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1012__A0  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0859__A1_N  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0856__B1  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0835__B2  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0827__A_N  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__D (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__C (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1067__A1  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1028__A1  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0832__A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0828__A_N  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__D (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__C (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._1028__A3  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0844__A_N  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0832__B1  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__C (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__D (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0842__A  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__C (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__C (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__D (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__C (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0898__A  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0893__B_N  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__C (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__D (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0921__A0  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0892__A  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0890__B  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__D (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__C (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__D (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0840__A_N  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0838__B_N  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__D (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__C (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0871__A2  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_AuI._0825__B2  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08840__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__C (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(net133));
 sky130_fd_sc_hd__fill_1 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1058 ();
endmodule

