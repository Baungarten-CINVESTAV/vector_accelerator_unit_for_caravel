VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Top_Module_4_ALU
  CLASS BLOCK ;
  FOREIGN Top_Module_4_ALU ;
  ORIGIN 0.000 0.000 ;
  SIZE 975.000 BY 1900.000 ;
  PIN ALU_Output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 1896.000 934.170 1899.000 ;
    END
  END ALU_Output[0]
  PIN ALU_Output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1336.240 4.000 1336.840 ;
    END
  END ALU_Output[100]
  PIN ALU_Output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 115.640 974.000 116.240 ;
    END
  END ALU_Output[101]
  PIN ALU_Output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1706.840 974.000 1707.440 ;
    END
  END ALU_Output[102]
  PIN ALU_Output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 1896.000 209.670 1899.000 ;
    END
  END ALU_Output[103]
  PIN ALU_Output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 581.440 974.000 582.040 ;
    END
  END ALU_Output[104]
  PIN ALU_Output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1686.440 974.000 1687.040 ;
    END
  END ALU_Output[105]
  PIN ALU_Output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 1896.000 592.850 1899.000 ;
    END
  END ALU_Output[106]
  PIN ALU_Output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1315.840 4.000 1316.440 ;
    END
  END ALU_Output[107]
  PIN ALU_Output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 221.040 974.000 221.640 ;
    END
  END ALU_Output[108]
  PIN ALU_Output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1040.440 4.000 1041.040 ;
    END
  END ALU_Output[109]
  PIN ALU_Output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 40.840 4.000 41.440 ;
    END
  END ALU_Output[10]
  PIN ALU_Output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 1896.000 573.530 1899.000 ;
    END
  END ALU_Output[110]
  PIN ALU_Output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1071.040 974.000 1071.640 ;
    END
  END ALU_Output[111]
  PIN ALU_Output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1485.840 4.000 1486.440 ;
    END
  END ALU_Output[112]
  PIN ALU_Output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1761.240 4.000 1761.840 ;
    END
  END ALU_Output[113]
  PIN ALU_Output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 306.040 974.000 306.640 ;
    END
  END ALU_Output[114]
  PIN ALU_Output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1145.840 4.000 1146.440 ;
    END
  END ALU_Output[115]
  PIN ALU_Output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 326.440 974.000 327.040 ;
    END
  END ALU_Output[116]
  PIN ALU_Output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 1.000 480.150 4.000 ;
    END
  END ALU_Output[117]
  PIN ALU_Output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 1896.000 654.030 1899.000 ;
    END
  END ALU_Output[118]
  PIN ALU_Output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 1.000 361.010 4.000 ;
    END
  END ALU_Output[119]
  PIN ALU_Output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 1896.000 270.850 1899.000 ;
    END
  END ALU_Output[11]
  PIN ALU_Output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1591.240 4.000 1591.840 ;
    END
  END ALU_Output[120]
  PIN ALU_Output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1295.440 4.000 1296.040 ;
    END
  END ALU_Output[121]
  PIN ALU_Output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1081.240 4.000 1081.840 ;
    END
  END ALU_Output[122]
  PIN ALU_Output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 486.240 4.000 486.840 ;
    END
  END ALU_Output[123]
  PIN ALU_Output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1281.840 974.000 1282.440 ;
    END
  END ALU_Output[124]
  PIN ALU_Output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 1896.000 251.530 1899.000 ;
    END
  END ALU_Output[125]
  PIN ALU_Output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 996.240 4.000 996.840 ;
    END
  END ALU_Output[126]
  PIN ALU_Output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 1.000 560.650 4.000 ;
    END
  END ALU_Output[127]
  PIN ALU_Output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1305.640 974.000 1306.240 ;
    END
  END ALU_Output[12]
  PIN ALU_Output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 1896.000 29.350 1899.000 ;
    END
  END ALU_Output[13]
  PIN ALU_Output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 411.440 974.000 412.040 ;
    END
  END ALU_Output[14]
  PIN ALU_Output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 71.440 974.000 72.040 ;
    END
  END ALU_Output[15]
  PIN ALU_Output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 1.000 583.190 4.000 ;
    END
  END ALU_Output[16]
  PIN ALU_Output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1230.840 4.000 1231.440 ;
    END
  END ALU_Output[17]
  PIN ALU_Output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1125.440 4.000 1126.040 ;
    END
  END ALU_Output[18]
  PIN ALU_Output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 156.440 974.000 157.040 ;
    END
  END ALU_Output[19]
  PIN ALU_Output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1781.640 4.000 1782.240 ;
    END
  END ALU_Output[1]
  PIN ALU_Output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 1.000 341.690 4.000 ;
    END
  END ALU_Output[20]
  PIN ALU_Output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 1896.000 550.990 1899.000 ;
    END
  END ALU_Output[21]
  PIN ALU_Output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 370.640 974.000 371.240 ;
    END
  END ALU_Output[22]
  PIN ALU_Output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 676.640 4.000 677.240 ;
    END
  END ALU_Output[23]
  PIN ALU_Output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 720.840 4.000 721.440 ;
    END
  END ALU_Output[24]
  PIN ALU_Output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 10.240 974.000 10.840 ;
    END
  END ALU_Output[25]
  PIN ALU_Output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 1896.000 67.990 1899.000 ;
    END
  END ALU_Output[26]
  PIN ALU_Output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 1.000 602.510 4.000 ;
    END
  END ALU_Output[27]
  PIN ALU_Output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 1896.000 470.490 1899.000 ;
    END
  END ALU_Output[28]
  PIN ALU_Output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1261.440 974.000 1262.040 ;
    END
  END ALU_Output[29]
  PIN ALU_Output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 1896.000 309.490 1899.000 ;
    END
  END ALU_Output[2]
  PIN ALU_Output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1887.040 4.000 1887.640 ;
    END
  END ALU_Output[30]
  PIN ALU_Output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1560.640 974.000 1561.240 ;
    END
  END ALU_Output[31]
  PIN ALU_Output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1740.840 4.000 1741.440 ;
    END
  END ALU_Output[32]
  PIN ALU_Output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 1.000 763.510 4.000 ;
    END
  END ALU_Output[33]
  PIN ALU_Output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 741.240 4.000 741.840 ;
    END
  END ALU_Output[34]
  PIN ALU_Output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1547.040 4.000 1547.640 ;
    END
  END ALU_Output[35]
  PIN ALU_Output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 1.000 77.650 4.000 ;
    END
  END ALU_Output[36]
  PIN ALU_Output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 846.640 4.000 847.240 ;
    END
  END ALU_Output[37]
  PIN ALU_Output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1451.840 974.000 1452.440 ;
    END
  END ALU_Output[38]
  PIN ALU_Output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 1.000 238.650 4.000 ;
    END
  END ALU_Output[39]
  PIN ALU_Output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1166.240 4.000 1166.840 ;
    END
  END ALU_Output[3]
  PIN ALU_Output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 496.440 974.000 497.040 ;
    END
  END ALU_Output[40]
  PIN ALU_Output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1791.840 974.000 1792.440 ;
    END
  END ALU_Output[41]
  PIN ALU_Output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 455.640 974.000 456.240 ;
    END
  END ALU_Output[42]
  PIN ALU_Output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 1.000 319.150 4.000 ;
    END
  END ALU_Output[43]
  PIN ALU_Output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1506.240 4.000 1506.840 ;
    END
  END ALU_Output[44]
  PIN ALU_Output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 265.240 974.000 265.840 ;
    END
  END ALU_Output[45]
  PIN ALU_Output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1866.640 4.000 1867.240 ;
    END
  END ALU_Output[46]
  PIN ALU_Output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 686.840 974.000 687.440 ;
    END
  END ALU_Output[47]
  PIN ALU_Output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 1896.000 370.670 1899.000 ;
    END
  END ALU_Output[48]
  PIN ALU_Output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 795.640 974.000 796.240 ;
    END
  END ALU_Output[49]
  PIN ALU_Output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 1896.000 109.850 1899.000 ;
    END
  END ALU_Output[4]
  PIN ALU_Output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1655.840 4.000 1656.440 ;
    END
  END ALU_Output[50]
  PIN ALU_Output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1676.240 4.000 1676.840 ;
    END
  END ALU_Output[51]
  PIN ALU_Output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 1896.000 834.350 1899.000 ;
    END
  END ALU_Output[52]
  PIN ALU_Output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 275.440 4.000 276.040 ;
    END
  END ALU_Output[53]
  PIN ALU_Output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 666.440 974.000 667.040 ;
    END
  END ALU_Output[54]
  PIN ALU_Output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1836.040 974.000 1836.640 ;
    END
  END ALU_Output[55]
  PIN ALU_Output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 1896.000 972.810 1899.000 ;
    END
  END ALU_Output[56]
  PIN ALU_Output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 1.000 158.150 4.000 ;
    END
  END ALU_Output[57]
  PIN ALU_Output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 1.000 702.330 4.000 ;
    END
  END ALU_Output[58]
  PIN ALU_Output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1876.840 974.000 1877.440 ;
    END
  END ALU_Output[59]
  PIN ALU_Output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 210.840 4.000 211.440 ;
    END
  END ALU_Output[5]
  PIN ALU_Output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1570.840 4.000 1571.440 ;
    END
  END ALU_Output[60]
  PIN ALU_Output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250 1896.000 895.530 1899.000 ;
    END
  END ALU_Output[61]
  PIN ALU_Output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 1.000 441.510 4.000 ;
    END
  END ALU_Output[62]
  PIN ALU_Output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 890.840 4.000 891.440 ;
    END
  END ALU_Output[63]
  PIN ALU_Output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 1.000 422.190 4.000 ;
    END
  END ALU_Output[64]
  PIN ALU_Output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 295.840 4.000 296.440 ;
    END
  END ALU_Output[65]
  PIN ALU_Output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 1896.000 171.030 1899.000 ;
    END
  END ALU_Output[66]
  PIN ALU_Output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1176.440 974.000 1177.040 ;
    END
  END ALU_Output[67]
  PIN ALU_Output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 625.640 974.000 626.240 ;
    END
  END ALU_Output[68]
  PIN ALU_Output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 1896.000 228.990 1899.000 ;
    END
  END ALU_Output[69]
  PIN ALU_Output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 1896.000 493.030 1899.000 ;
    END
  END ALU_Output[6]
  PIN ALU_Output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 1.000 219.330 4.000 ;
    END
  END ALU_Output[70]
  PIN ALU_Output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1326.040 974.000 1326.640 ;
    END
  END ALU_Output[71]
  PIN ALU_Output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1462.040 4.000 1462.640 ;
    END
  END ALU_Output[72]
  PIN ALU_Output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 136.040 974.000 136.640 ;
    END
  END ALU_Output[73]
  PIN ALU_Output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 1896.000 734.530 1899.000 ;
    END
  END ALU_Output[74]
  PIN ALU_Output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 1.000 541.330 4.000 ;
    END
  END ALU_Output[75]
  PIN ALU_Output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 350.240 974.000 350.840 ;
    END
  END ALU_Output[76]
  PIN ALU_Output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 1896.000 631.490 1899.000 ;
    END
  END ALU_Output[77]
  PIN ALU_Output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 561.040 974.000 561.640 ;
    END
  END ALU_Output[78]
  PIN ALU_Output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 826.240 4.000 826.840 ;
    END
  END ALU_Output[79]
  PIN ALU_Output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1271.640 4.000 1272.240 ;
    END
  END ALU_Output[7]
  PIN ALU_Output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 1896.000 914.850 1899.000 ;
    END
  END ALU_Output[80]
  PIN ALU_Output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1825.840 4.000 1826.440 ;
    END
  END ALU_Output[81]
  PIN ALU_Output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 550.840 4.000 551.440 ;
    END
  END ALU_Output[82]
  PIN ALU_Output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1802.040 4.000 1802.640 ;
    END
  END ALU_Output[83]
  PIN ALU_Output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1896.000 48.670 1899.000 ;
    END
  END ALU_Output[84]
  PIN ALU_Output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 1896.000 129.170 1899.000 ;
    END
  END ALU_Output[85]
  PIN ALU_Output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 81.640 4.000 82.240 ;
    END
  END ALU_Output[86]
  PIN ALU_Output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 476.040 974.000 476.640 ;
    END
  END ALU_Output[87]
  PIN ALU_Output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1026.840 974.000 1027.440 ;
    END
  END ALU_Output[88]
  PIN ALU_Output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 421.640 4.000 422.240 ;
    END
  END ALU_Output[89]
  PIN ALU_Output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1241.040 974.000 1241.640 ;
    END
  END ALU_Output[8]
  PIN ALU_Output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 125.840 4.000 126.440 ;
    END
  END ALU_Output[90]
  PIN ALU_Output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1846.240 4.000 1846.840 ;
    END
  END ALU_Output[91]
  PIN ALU_Output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 1.000 863.330 4.000 ;
    END
  END ALU_Output[92]
  PIN ALU_Output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1346.440 974.000 1347.040 ;
    END
  END ALU_Output[93]
  PIN ALU_Output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 1.000 180.690 4.000 ;
    END
  END ALU_Output[94]
  PIN ALU_Output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 700.440 4.000 701.040 ;
    END
  END ALU_Output[95]
  PIN ALU_Output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1356.640 4.000 1357.240 ;
    END
  END ALU_Output[96]
  PIN ALU_Output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 1896.000 148.490 1899.000 ;
    END
  END ALU_Output[97]
  PIN ALU_Output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 901.040 974.000 901.640 ;
    END
  END ALU_Output[98]
  PIN ALU_Output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1666.040 974.000 1666.640 ;
    END
  END ALU_Output[99]
  PIN ALU_Output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 880.640 974.000 881.240 ;
    END
  END ALU_Output[9]
  PIN Exception[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 1.000 502.690 4.000 ;
    END
  END Exception[0]
  PIN Exception[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1220.640 974.000 1221.240 ;
    END
  END Exception[1]
  PIN Exception[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 761.640 4.000 762.240 ;
    END
  END Exception[2]
  PIN Exception[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 591.640 4.000 592.240 ;
    END
  END Exception[3]
  PIN Operation[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 1.000 782.830 4.000 ;
    END
  END Operation[0]
  PIN Operation[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 251.640 4.000 252.240 ;
    END
  END Operation[1]
  PIN Operation[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 1896.000 753.850 1899.000 ;
    END
  END Operation[2]
  PIN Operation[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1196.840 974.000 1197.440 ;
    END
  END Operation[3]
  PIN Overflow[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 200.640 974.000 201.240 ;
    END
  END Overflow[0]
  PIN Overflow[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 530.440 4.000 531.040 ;
    END
  END Overflow[1]
  PIN Overflow[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1400.840 4.000 1401.440 ;
    END
  END Overflow[2]
  PIN Overflow[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1186.640 4.000 1187.240 ;
    END
  END Overflow[3]
  PIN Underflow[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1717.040 4.000 1717.640 ;
    END
  END Underflow[0]
  PIN Underflow[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1366.840 974.000 1367.440 ;
    END
  END Underflow[1]
  PIN Underflow[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 1.000 844.010 4.000 ;
    END
  END Underflow[2]
  PIN Underflow[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 316.240 4.000 316.840 ;
    END
  END Underflow[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 1.000 802.150 4.000 ;
    END
  END clk
  PIN iCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1526.640 4.000 1527.240 ;
    END
  END iCE
  PIN i_operand_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 856.840 974.000 857.440 ;
    END
  END i_operand_sel
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 1896.000 431.850 1899.000 ;
    END
  END i_rst
  PIN operand[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 1896.000 872.990 1899.000 ;
    END
  END operand[0]
  PIN operand[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1896.000 451.170 1899.000 ;
    END
  END operand[100]
  PIN operand[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 836.440 974.000 837.040 ;
    END
  END operand[101]
  PIN operand[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1621.840 974.000 1622.440 ;
    END
  END operand[102]
  PIN operand[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 710.640 974.000 711.240 ;
    END
  END operand[103]
  PIN operand[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 231.240 4.000 231.840 ;
    END
  END operand[104]
  PIN operand[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1411.040 974.000 1411.640 ;
    END
  END operand[105]
  PIN operand[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 241.440 974.000 242.040 ;
    END
  END operand[106]
  PIN operand[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1771.440 974.000 1772.040 ;
    END
  END operand[107]
  PIN operand[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 51.040 974.000 51.640 ;
    END
  END operand[108]
  PIN operand[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 1896.000 351.350 1899.000 ;
    END
  END operand[109]
  PIN operand[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 1.000 138.830 4.000 ;
    END
  END operand[10]
  PIN operand[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 731.040 974.000 731.640 ;
    END
  END operand[110]
  PIN operand[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 1.000 621.830 4.000 ;
    END
  END operand[111]
  PIN operand[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 921.440 974.000 922.040 ;
    END
  END operand[112]
  PIN operand[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 465.840 4.000 466.440 ;
    END
  END operand[113]
  PIN operand[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1016.640 4.000 1017.240 ;
    END
  END operand[114]
  PIN operand[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 1896.000 673.350 1899.000 ;
    END
  END operand[115]
  PIN operand[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1536.840 974.000 1537.440 ;
    END
  END operand[116]
  PIN operand[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1091.440 974.000 1092.040 ;
    END
  END operand[117]
  PIN operand[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 360.440 4.000 361.040 ;
    END
  END operand[118]
  PIN operand[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 1896.000 692.670 1899.000 ;
    END
  END operand[119]
  PIN operand[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 955.440 4.000 956.040 ;
    END
  END operand[11]
  PIN operand[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 146.240 4.000 146.840 ;
    END
  END operand[120]
  PIN operand[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 506.640 4.000 507.240 ;
    END
  END operand[121]
  PIN operand[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1441.640 4.000 1442.240 ;
    END
  END operand[122]
  PIN operand[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 1896.000 792.490 1899.000 ;
    END
  END operand[123]
  PIN operand[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 1896.000 332.030 1899.000 ;
    END
  END operand[124]
  PIN operand[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 805.840 4.000 806.440 ;
    END
  END operand[125]
  PIN operand[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 911.240 4.000 911.840 ;
    END
  END operand[126]
  PIN operand[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1111.840 974.000 1112.440 ;
    END
  END operand[127]
  PIN operand[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1050.640 974.000 1051.240 ;
    END
  END operand[12]
  PIN operand[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 380.840 4.000 381.440 ;
    END
  END operand[13]
  PIN operand[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 965.640 974.000 966.240 ;
    END
  END operand[14]
  PIN operand[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 601.840 974.000 602.440 ;
    END
  END operand[15]
  PIN operand[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 180.240 974.000 180.840 ;
    END
  END operand[16]
  PIN operand[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 975.840 4.000 976.440 ;
    END
  END operand[17]
  PIN operand[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1581.040 974.000 1581.640 ;
    END
  END operand[18]
  PIN operand[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 1.000 683.010 4.000 ;
    END
  END operand[19]
  PIN operand[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 1.000 963.150 4.000 ;
    END
  END operand[1]
  PIN operand[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 516.840 974.000 517.440 ;
    END
  END operand[20]
  PIN operand[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1896.000 290.170 1899.000 ;
    END
  END operand[21]
  PIN operand[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 1.000 663.690 4.000 ;
    END
  END operand[22]
  PIN operand[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 1.000 119.510 4.000 ;
    END
  END operand[23]
  PIN operand[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 166.640 4.000 167.240 ;
    END
  END operand[24]
  PIN operand[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1006.440 974.000 1007.040 ;
    END
  END operand[25]
  PIN operand[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1475.640 974.000 1476.240 ;
    END
  END operand[26]
  PIN operand[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 1.000 460.830 4.000 ;
    END
  END operand[27]
  PIN operand[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1815.640 974.000 1816.240 ;
    END
  END operand[28]
  PIN operand[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 61.240 4.000 61.840 ;
    END
  END operand[29]
  PIN operand[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 1.000 943.830 4.000 ;
    END
  END operand[2]
  PIN operand[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1856.440 974.000 1857.040 ;
    END
  END operand[30]
  PIN operand[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 1.000 924.510 4.000 ;
    END
  END operand[31]
  PIN operand[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 1.000 380.330 4.000 ;
    END
  END operand[32]
  PIN operand[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 1.000 58.330 4.000 ;
    END
  END operand[33]
  PIN operand[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 285.640 974.000 286.240 ;
    END
  END operand[34]
  PIN operand[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 646.040 974.000 646.640 ;
    END
  END operand[35]
  PIN operand[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 1896.000 412.530 1899.000 ;
    END
  END operand[36]
  PIN operand[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1431.440 974.000 1432.040 ;
    END
  END operand[37]
  PIN operand[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1611.640 4.000 1612.240 ;
    END
  END operand[38]
  PIN operand[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1696.640 4.000 1697.240 ;
    END
  END operand[39]
  PIN operand[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 105.440 4.000 106.040 ;
    END
  END operand[3]
  PIN operand[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 1.000 39.010 4.000 ;
    END
  END operand[40]
  PIN operand[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 1.000 261.190 4.000 ;
    END
  END operand[41]
  PIN operand[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 986.040 974.000 986.640 ;
    END
  END operand[42]
  PIN operand[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1.000 721.650 4.000 ;
    END
  END operand[43]
  PIN operand[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 1896.000 815.030 1899.000 ;
    END
  END operand[44]
  PIN operand[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1751.040 974.000 1751.640 ;
    END
  END operand[45]
  PIN operand[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 1896.000 10.030 1899.000 ;
    END
  END operand[46]
  PIN operand[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 931.640 4.000 932.240 ;
    END
  END operand[47]
  PIN operand[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1135.640 974.000 1136.240 ;
    END
  END operand[48]
  PIN operand[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1730.640 974.000 1731.240 ;
    END
  END operand[49]
  PIN operand[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1251.240 4.000 1251.840 ;
    END
  END operand[4]
  PIN operand[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1390.640 974.000 1391.240 ;
    END
  END operand[50]
  PIN operand[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 771.840 974.000 772.440 ;
    END
  END operand[51]
  PIN operand[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 1.000 882.650 4.000 ;
    END
  END operand[52]
  PIN operand[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 1896.000 953.490 1899.000 ;
    END
  END operand[53]
  PIN operand[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 1896.000 190.350 1899.000 ;
    END
  END operand[54]
  PIN operand[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 1.000 399.650 4.000 ;
    END
  END operand[55]
  PIN operand[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 785.440 4.000 786.040 ;
    END
  END operand[56]
  PIN operand[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 571.240 4.000 571.840 ;
    END
  END operand[57]
  PIN operand[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 751.440 974.000 752.040 ;
    END
  END operand[58]
  PIN operand[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1101.640 4.000 1102.240 ;
    END
  END operand[59]
  PIN operand[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 391.040 974.000 391.640 ;
    END
  END operand[5]
  PIN operand[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 1.000 200.010 4.000 ;
    END
  END operand[60]
  PIN operand[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 1.000 641.150 4.000 ;
    END
  END operand[61]
  PIN operand[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 941.840 974.000 942.440 ;
    END
  END operand[62]
  PIN operand[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1896.000 853.670 1899.000 ;
    END
  END operand[63]
  PIN operand[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1601.440 974.000 1602.040 ;
    END
  END operand[64]
  PIN operand[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 435.240 974.000 435.840 ;
    END
  END operand[65]
  PIN operand[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 445.440 4.000 446.040 ;
    END
  END operand[66]
  PIN operand[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 20.440 4.000 21.040 ;
    END
  END operand[67]
  PIN operand[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 1.000 19.690 4.000 ;
    END
  END operand[68]
  PIN operand[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1645.640 974.000 1646.240 ;
    END
  END operand[69]
  PIN operand[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 1896.000 773.170 1899.000 ;
    END
  END operand[6]
  PIN operand[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 540.640 974.000 541.240 ;
    END
  END operand[70]
  PIN operand[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 1896.000 711.990 1899.000 ;
    END
  END operand[71]
  PIN operand[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 615.440 4.000 616.040 ;
    END
  END operand[72]
  PIN operand[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 656.240 4.000 656.840 ;
    END
  END operand[73]
  PIN operand[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.910 1.000 905.190 4.000 ;
    END
  END operand[74]
  PIN operand[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 1.000 0.370 4.000 ;
    END
  END operand[75]
  PIN operand[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 95.240 974.000 95.840 ;
    END
  END operand[76]
  PIN operand[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 870.440 4.000 871.040 ;
    END
  END operand[77]
  PIN operand[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1421.240 4.000 1421.840 ;
    END
  END operand[78]
  PIN operand[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 401.240 4.000 401.840 ;
    END
  END operand[79]
  PIN operand[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 635.840 4.000 636.440 ;
    END
  END operand[7]
  PIN operand[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 1.000 280.510 4.000 ;
    END
  END operand[80]
  PIN operand[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 1.000 100.190 4.000 ;
    END
  END operand[81]
  PIN operand[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 1896.000 389.990 1899.000 ;
    END
  END operand[82]
  PIN operand[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 1896.000 90.530 1899.000 ;
    END
  END operand[83]
  PIN operand[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 1.000 744.190 4.000 ;
    END
  END operand[84]
  PIN operand[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1896.000 612.170 1899.000 ;
    END
  END operand[85]
  PIN operand[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 816.040 974.000 816.640 ;
    END
  END operand[86]
  PIN operand[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1060.840 4.000 1061.440 ;
    END
  END operand[87]
  PIN operand[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1516.440 974.000 1517.040 ;
    END
  END operand[88]
  PIN operand[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 1.000 299.830 4.000 ;
    END
  END operand[89]
  PIN operand[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 1.000 522.010 4.000 ;
    END
  END operand[8]
  PIN operand[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 190.440 4.000 191.040 ;
    END
  END operand[90]
  PIN operand[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1496.040 974.000 1496.640 ;
    END
  END operand[91]
  PIN operand[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 1.000 824.690 4.000 ;
    END
  END operand[92]
  PIN operand[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 1896.000 531.670 1899.000 ;
    END
  END operand[93]
  PIN operand[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 1896.000 512.350 1899.000 ;
    END
  END operand[94]
  PIN operand[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1380.440 4.000 1381.040 ;
    END
  END operand[95]
  PIN operand[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1632.040 4.000 1632.640 ;
    END
  END operand[96]
  PIN operand[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 30.640 974.000 31.240 ;
    END
  END operand[97]
  PIN operand[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 336.640 4.000 337.240 ;
    END
  END operand[98]
  PIN operand[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.000 1210.440 4.000 1211.040 ;
    END
  END operand[99]
  PIN operand[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 971.000 1156.040 974.000 1156.640 ;
    END
  END operand[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1887.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1887.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1887.920 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 969.220 1887.765 ;
      LAYER met1 ;
        RECT 0.070 10.640 974.670 1887.920 ;
      LAYER met2 ;
        RECT 0.100 1895.720 9.470 1896.000 ;
        RECT 10.310 1895.720 28.790 1896.000 ;
        RECT 29.630 1895.720 48.110 1896.000 ;
        RECT 48.950 1895.720 67.430 1896.000 ;
        RECT 68.270 1895.720 89.970 1896.000 ;
        RECT 90.810 1895.720 109.290 1896.000 ;
        RECT 110.130 1895.720 128.610 1896.000 ;
        RECT 129.450 1895.720 147.930 1896.000 ;
        RECT 148.770 1895.720 170.470 1896.000 ;
        RECT 171.310 1895.720 189.790 1896.000 ;
        RECT 190.630 1895.720 209.110 1896.000 ;
        RECT 209.950 1895.720 228.430 1896.000 ;
        RECT 229.270 1895.720 250.970 1896.000 ;
        RECT 251.810 1895.720 270.290 1896.000 ;
        RECT 271.130 1895.720 289.610 1896.000 ;
        RECT 290.450 1895.720 308.930 1896.000 ;
        RECT 309.770 1895.720 331.470 1896.000 ;
        RECT 332.310 1895.720 350.790 1896.000 ;
        RECT 351.630 1895.720 370.110 1896.000 ;
        RECT 370.950 1895.720 389.430 1896.000 ;
        RECT 390.270 1895.720 411.970 1896.000 ;
        RECT 412.810 1895.720 431.290 1896.000 ;
        RECT 432.130 1895.720 450.610 1896.000 ;
        RECT 451.450 1895.720 469.930 1896.000 ;
        RECT 470.770 1895.720 492.470 1896.000 ;
        RECT 493.310 1895.720 511.790 1896.000 ;
        RECT 512.630 1895.720 531.110 1896.000 ;
        RECT 531.950 1895.720 550.430 1896.000 ;
        RECT 551.270 1895.720 572.970 1896.000 ;
        RECT 573.810 1895.720 592.290 1896.000 ;
        RECT 593.130 1895.720 611.610 1896.000 ;
        RECT 612.450 1895.720 630.930 1896.000 ;
        RECT 631.770 1895.720 653.470 1896.000 ;
        RECT 654.310 1895.720 672.790 1896.000 ;
        RECT 673.630 1895.720 692.110 1896.000 ;
        RECT 692.950 1895.720 711.430 1896.000 ;
        RECT 712.270 1895.720 733.970 1896.000 ;
        RECT 734.810 1895.720 753.290 1896.000 ;
        RECT 754.130 1895.720 772.610 1896.000 ;
        RECT 773.450 1895.720 791.930 1896.000 ;
        RECT 792.770 1895.720 814.470 1896.000 ;
        RECT 815.310 1895.720 833.790 1896.000 ;
        RECT 834.630 1895.720 853.110 1896.000 ;
        RECT 853.950 1895.720 872.430 1896.000 ;
        RECT 873.270 1895.720 894.970 1896.000 ;
        RECT 895.810 1895.720 914.290 1896.000 ;
        RECT 915.130 1895.720 933.610 1896.000 ;
        RECT 934.450 1895.720 952.930 1896.000 ;
        RECT 953.770 1895.720 972.250 1896.000 ;
        RECT 973.090 1895.720 974.650 1896.000 ;
        RECT 0.100 4.280 974.650 1895.720 ;
        RECT 0.650 3.670 19.130 4.280 ;
        RECT 19.970 3.670 38.450 4.280 ;
        RECT 39.290 3.670 57.770 4.280 ;
        RECT 58.610 3.670 77.090 4.280 ;
        RECT 77.930 3.670 99.630 4.280 ;
        RECT 100.470 3.670 118.950 4.280 ;
        RECT 119.790 3.670 138.270 4.280 ;
        RECT 139.110 3.670 157.590 4.280 ;
        RECT 158.430 3.670 180.130 4.280 ;
        RECT 180.970 3.670 199.450 4.280 ;
        RECT 200.290 3.670 218.770 4.280 ;
        RECT 219.610 3.670 238.090 4.280 ;
        RECT 238.930 3.670 260.630 4.280 ;
        RECT 261.470 3.670 279.950 4.280 ;
        RECT 280.790 3.670 299.270 4.280 ;
        RECT 300.110 3.670 318.590 4.280 ;
        RECT 319.430 3.670 341.130 4.280 ;
        RECT 341.970 3.670 360.450 4.280 ;
        RECT 361.290 3.670 379.770 4.280 ;
        RECT 380.610 3.670 399.090 4.280 ;
        RECT 399.930 3.670 421.630 4.280 ;
        RECT 422.470 3.670 440.950 4.280 ;
        RECT 441.790 3.670 460.270 4.280 ;
        RECT 461.110 3.670 479.590 4.280 ;
        RECT 480.430 3.670 502.130 4.280 ;
        RECT 502.970 3.670 521.450 4.280 ;
        RECT 522.290 3.670 540.770 4.280 ;
        RECT 541.610 3.670 560.090 4.280 ;
        RECT 560.930 3.670 582.630 4.280 ;
        RECT 583.470 3.670 601.950 4.280 ;
        RECT 602.790 3.670 621.270 4.280 ;
        RECT 622.110 3.670 640.590 4.280 ;
        RECT 641.430 3.670 663.130 4.280 ;
        RECT 663.970 3.670 682.450 4.280 ;
        RECT 683.290 3.670 701.770 4.280 ;
        RECT 702.610 3.670 721.090 4.280 ;
        RECT 721.930 3.670 743.630 4.280 ;
        RECT 744.470 3.670 762.950 4.280 ;
        RECT 763.790 3.670 782.270 4.280 ;
        RECT 783.110 3.670 801.590 4.280 ;
        RECT 802.430 3.670 824.130 4.280 ;
        RECT 824.970 3.670 843.450 4.280 ;
        RECT 844.290 3.670 862.770 4.280 ;
        RECT 863.610 3.670 882.090 4.280 ;
        RECT 882.930 3.670 904.630 4.280 ;
        RECT 905.470 3.670 923.950 4.280 ;
        RECT 924.790 3.670 943.270 4.280 ;
        RECT 944.110 3.670 962.590 4.280 ;
        RECT 963.430 3.670 974.650 4.280 ;
      LAYER met3 ;
        RECT 4.400 1886.640 974.890 1887.845 ;
        RECT 4.000 1877.840 974.890 1886.640 ;
        RECT 4.000 1876.440 970.600 1877.840 ;
        RECT 974.400 1876.440 974.890 1877.840 ;
        RECT 4.000 1867.640 974.890 1876.440 ;
        RECT 4.400 1866.240 974.890 1867.640 ;
        RECT 4.000 1857.440 974.890 1866.240 ;
        RECT 4.000 1856.040 970.600 1857.440 ;
        RECT 974.400 1856.040 974.890 1857.440 ;
        RECT 4.000 1847.240 974.890 1856.040 ;
        RECT 4.400 1845.840 974.890 1847.240 ;
        RECT 4.000 1837.040 974.890 1845.840 ;
        RECT 4.000 1835.640 970.600 1837.040 ;
        RECT 974.400 1835.640 974.890 1837.040 ;
        RECT 4.000 1826.840 974.890 1835.640 ;
        RECT 4.400 1825.440 974.890 1826.840 ;
        RECT 4.000 1816.640 974.890 1825.440 ;
        RECT 4.000 1815.240 970.600 1816.640 ;
        RECT 974.400 1815.240 974.890 1816.640 ;
        RECT 4.000 1803.040 974.890 1815.240 ;
        RECT 4.400 1801.640 974.890 1803.040 ;
        RECT 4.000 1792.840 974.890 1801.640 ;
        RECT 4.000 1791.440 970.600 1792.840 ;
        RECT 974.400 1791.440 974.890 1792.840 ;
        RECT 4.000 1782.640 974.890 1791.440 ;
        RECT 4.400 1781.240 974.890 1782.640 ;
        RECT 4.000 1772.440 974.890 1781.240 ;
        RECT 4.000 1771.040 970.600 1772.440 ;
        RECT 974.400 1771.040 974.890 1772.440 ;
        RECT 4.000 1762.240 974.890 1771.040 ;
        RECT 4.400 1760.840 974.890 1762.240 ;
        RECT 4.000 1752.040 974.890 1760.840 ;
        RECT 4.000 1750.640 970.600 1752.040 ;
        RECT 974.400 1750.640 974.890 1752.040 ;
        RECT 4.000 1741.840 974.890 1750.640 ;
        RECT 4.400 1740.440 974.890 1741.840 ;
        RECT 4.000 1731.640 974.890 1740.440 ;
        RECT 4.000 1730.240 970.600 1731.640 ;
        RECT 974.400 1730.240 974.890 1731.640 ;
        RECT 4.000 1718.040 974.890 1730.240 ;
        RECT 4.400 1716.640 974.890 1718.040 ;
        RECT 4.000 1707.840 974.890 1716.640 ;
        RECT 4.000 1706.440 970.600 1707.840 ;
        RECT 974.400 1706.440 974.890 1707.840 ;
        RECT 4.000 1697.640 974.890 1706.440 ;
        RECT 4.400 1696.240 974.890 1697.640 ;
        RECT 4.000 1687.440 974.890 1696.240 ;
        RECT 4.000 1686.040 970.600 1687.440 ;
        RECT 974.400 1686.040 974.890 1687.440 ;
        RECT 4.000 1677.240 974.890 1686.040 ;
        RECT 4.400 1675.840 974.890 1677.240 ;
        RECT 4.000 1667.040 974.890 1675.840 ;
        RECT 4.000 1665.640 970.600 1667.040 ;
        RECT 974.400 1665.640 974.890 1667.040 ;
        RECT 4.000 1656.840 974.890 1665.640 ;
        RECT 4.400 1655.440 974.890 1656.840 ;
        RECT 4.000 1646.640 974.890 1655.440 ;
        RECT 4.000 1645.240 970.600 1646.640 ;
        RECT 974.400 1645.240 974.890 1646.640 ;
        RECT 4.000 1633.040 974.890 1645.240 ;
        RECT 4.400 1631.640 974.890 1633.040 ;
        RECT 4.000 1622.840 974.890 1631.640 ;
        RECT 4.000 1621.440 970.600 1622.840 ;
        RECT 974.400 1621.440 974.890 1622.840 ;
        RECT 4.000 1612.640 974.890 1621.440 ;
        RECT 4.400 1611.240 974.890 1612.640 ;
        RECT 4.000 1602.440 974.890 1611.240 ;
        RECT 4.000 1601.040 970.600 1602.440 ;
        RECT 974.400 1601.040 974.890 1602.440 ;
        RECT 4.000 1592.240 974.890 1601.040 ;
        RECT 4.400 1590.840 974.890 1592.240 ;
        RECT 4.000 1582.040 974.890 1590.840 ;
        RECT 4.000 1580.640 970.600 1582.040 ;
        RECT 974.400 1580.640 974.890 1582.040 ;
        RECT 4.000 1571.840 974.890 1580.640 ;
        RECT 4.400 1570.440 974.890 1571.840 ;
        RECT 4.000 1561.640 974.890 1570.440 ;
        RECT 4.000 1560.240 970.600 1561.640 ;
        RECT 974.400 1560.240 974.890 1561.640 ;
        RECT 4.000 1548.040 974.890 1560.240 ;
        RECT 4.400 1546.640 974.890 1548.040 ;
        RECT 4.000 1537.840 974.890 1546.640 ;
        RECT 4.000 1536.440 970.600 1537.840 ;
        RECT 974.400 1536.440 974.890 1537.840 ;
        RECT 4.000 1527.640 974.890 1536.440 ;
        RECT 4.400 1526.240 974.890 1527.640 ;
        RECT 4.000 1517.440 974.890 1526.240 ;
        RECT 4.000 1516.040 970.600 1517.440 ;
        RECT 974.400 1516.040 974.890 1517.440 ;
        RECT 4.000 1507.240 974.890 1516.040 ;
        RECT 4.400 1505.840 974.890 1507.240 ;
        RECT 4.000 1497.040 974.890 1505.840 ;
        RECT 4.000 1495.640 970.600 1497.040 ;
        RECT 974.400 1495.640 974.890 1497.040 ;
        RECT 4.000 1486.840 974.890 1495.640 ;
        RECT 4.400 1485.440 974.890 1486.840 ;
        RECT 4.000 1476.640 974.890 1485.440 ;
        RECT 4.000 1475.240 970.600 1476.640 ;
        RECT 974.400 1475.240 974.890 1476.640 ;
        RECT 4.000 1463.040 974.890 1475.240 ;
        RECT 4.400 1461.640 974.890 1463.040 ;
        RECT 4.000 1452.840 974.890 1461.640 ;
        RECT 4.000 1451.440 970.600 1452.840 ;
        RECT 974.400 1451.440 974.890 1452.840 ;
        RECT 4.000 1442.640 974.890 1451.440 ;
        RECT 4.400 1441.240 974.890 1442.640 ;
        RECT 4.000 1432.440 974.890 1441.240 ;
        RECT 4.000 1431.040 970.600 1432.440 ;
        RECT 974.400 1431.040 974.890 1432.440 ;
        RECT 4.000 1422.240 974.890 1431.040 ;
        RECT 4.400 1420.840 974.890 1422.240 ;
        RECT 4.000 1412.040 974.890 1420.840 ;
        RECT 4.000 1410.640 970.600 1412.040 ;
        RECT 974.400 1410.640 974.890 1412.040 ;
        RECT 4.000 1401.840 974.890 1410.640 ;
        RECT 4.400 1400.440 974.890 1401.840 ;
        RECT 4.000 1391.640 974.890 1400.440 ;
        RECT 4.000 1390.240 970.600 1391.640 ;
        RECT 974.400 1390.240 974.890 1391.640 ;
        RECT 4.000 1381.440 974.890 1390.240 ;
        RECT 4.400 1380.040 974.890 1381.440 ;
        RECT 4.000 1367.840 974.890 1380.040 ;
        RECT 4.000 1366.440 970.600 1367.840 ;
        RECT 974.400 1366.440 974.890 1367.840 ;
        RECT 4.000 1357.640 974.890 1366.440 ;
        RECT 4.400 1356.240 974.890 1357.640 ;
        RECT 4.000 1347.440 974.890 1356.240 ;
        RECT 4.000 1346.040 970.600 1347.440 ;
        RECT 974.400 1346.040 974.890 1347.440 ;
        RECT 4.000 1337.240 974.890 1346.040 ;
        RECT 4.400 1335.840 974.890 1337.240 ;
        RECT 4.000 1327.040 974.890 1335.840 ;
        RECT 4.000 1325.640 970.600 1327.040 ;
        RECT 974.400 1325.640 974.890 1327.040 ;
        RECT 4.000 1316.840 974.890 1325.640 ;
        RECT 4.400 1315.440 974.890 1316.840 ;
        RECT 4.000 1306.640 974.890 1315.440 ;
        RECT 4.000 1305.240 970.600 1306.640 ;
        RECT 974.400 1305.240 974.890 1306.640 ;
        RECT 4.000 1296.440 974.890 1305.240 ;
        RECT 4.400 1295.040 974.890 1296.440 ;
        RECT 4.000 1282.840 974.890 1295.040 ;
        RECT 4.000 1281.440 970.600 1282.840 ;
        RECT 974.400 1281.440 974.890 1282.840 ;
        RECT 4.000 1272.640 974.890 1281.440 ;
        RECT 4.400 1271.240 974.890 1272.640 ;
        RECT 4.000 1262.440 974.890 1271.240 ;
        RECT 4.000 1261.040 970.600 1262.440 ;
        RECT 974.400 1261.040 974.890 1262.440 ;
        RECT 4.000 1252.240 974.890 1261.040 ;
        RECT 4.400 1250.840 974.890 1252.240 ;
        RECT 4.000 1242.040 974.890 1250.840 ;
        RECT 4.000 1240.640 970.600 1242.040 ;
        RECT 974.400 1240.640 974.890 1242.040 ;
        RECT 4.000 1231.840 974.890 1240.640 ;
        RECT 4.400 1230.440 974.890 1231.840 ;
        RECT 4.000 1221.640 974.890 1230.440 ;
        RECT 4.000 1220.240 970.600 1221.640 ;
        RECT 974.400 1220.240 974.890 1221.640 ;
        RECT 4.000 1211.440 974.890 1220.240 ;
        RECT 4.400 1210.040 974.890 1211.440 ;
        RECT 4.000 1197.840 974.890 1210.040 ;
        RECT 4.000 1196.440 970.600 1197.840 ;
        RECT 974.400 1196.440 974.890 1197.840 ;
        RECT 4.000 1187.640 974.890 1196.440 ;
        RECT 4.400 1186.240 974.890 1187.640 ;
        RECT 4.000 1177.440 974.890 1186.240 ;
        RECT 4.000 1176.040 970.600 1177.440 ;
        RECT 974.400 1176.040 974.890 1177.440 ;
        RECT 4.000 1167.240 974.890 1176.040 ;
        RECT 4.400 1165.840 974.890 1167.240 ;
        RECT 4.000 1157.040 974.890 1165.840 ;
        RECT 4.000 1155.640 970.600 1157.040 ;
        RECT 974.400 1155.640 974.890 1157.040 ;
        RECT 4.000 1146.840 974.890 1155.640 ;
        RECT 4.400 1145.440 974.890 1146.840 ;
        RECT 4.000 1136.640 974.890 1145.440 ;
        RECT 4.000 1135.240 970.600 1136.640 ;
        RECT 974.400 1135.240 974.890 1136.640 ;
        RECT 4.000 1126.440 974.890 1135.240 ;
        RECT 4.400 1125.040 974.890 1126.440 ;
        RECT 4.000 1112.840 974.890 1125.040 ;
        RECT 4.000 1111.440 970.600 1112.840 ;
        RECT 974.400 1111.440 974.890 1112.840 ;
        RECT 4.000 1102.640 974.890 1111.440 ;
        RECT 4.400 1101.240 974.890 1102.640 ;
        RECT 4.000 1092.440 974.890 1101.240 ;
        RECT 4.000 1091.040 970.600 1092.440 ;
        RECT 974.400 1091.040 974.890 1092.440 ;
        RECT 4.000 1082.240 974.890 1091.040 ;
        RECT 4.400 1080.840 974.890 1082.240 ;
        RECT 4.000 1072.040 974.890 1080.840 ;
        RECT 4.000 1070.640 970.600 1072.040 ;
        RECT 974.400 1070.640 974.890 1072.040 ;
        RECT 4.000 1061.840 974.890 1070.640 ;
        RECT 4.400 1060.440 974.890 1061.840 ;
        RECT 4.000 1051.640 974.890 1060.440 ;
        RECT 4.000 1050.240 970.600 1051.640 ;
        RECT 974.400 1050.240 974.890 1051.640 ;
        RECT 4.000 1041.440 974.890 1050.240 ;
        RECT 4.400 1040.040 974.890 1041.440 ;
        RECT 4.000 1027.840 974.890 1040.040 ;
        RECT 4.000 1026.440 970.600 1027.840 ;
        RECT 974.400 1026.440 974.890 1027.840 ;
        RECT 4.000 1017.640 974.890 1026.440 ;
        RECT 4.400 1016.240 974.890 1017.640 ;
        RECT 4.000 1007.440 974.890 1016.240 ;
        RECT 4.000 1006.040 970.600 1007.440 ;
        RECT 974.400 1006.040 974.890 1007.440 ;
        RECT 4.000 997.240 974.890 1006.040 ;
        RECT 4.400 995.840 974.890 997.240 ;
        RECT 4.000 987.040 974.890 995.840 ;
        RECT 4.000 985.640 970.600 987.040 ;
        RECT 974.400 985.640 974.890 987.040 ;
        RECT 4.000 976.840 974.890 985.640 ;
        RECT 4.400 975.440 974.890 976.840 ;
        RECT 4.000 966.640 974.890 975.440 ;
        RECT 4.000 965.240 970.600 966.640 ;
        RECT 974.400 965.240 974.890 966.640 ;
        RECT 4.000 956.440 974.890 965.240 ;
        RECT 4.400 955.040 974.890 956.440 ;
        RECT 4.000 942.840 974.890 955.040 ;
        RECT 4.000 941.440 970.600 942.840 ;
        RECT 974.400 941.440 974.890 942.840 ;
        RECT 4.000 932.640 974.890 941.440 ;
        RECT 4.400 931.240 974.890 932.640 ;
        RECT 4.000 922.440 974.890 931.240 ;
        RECT 4.000 921.040 970.600 922.440 ;
        RECT 974.400 921.040 974.890 922.440 ;
        RECT 4.000 912.240 974.890 921.040 ;
        RECT 4.400 910.840 974.890 912.240 ;
        RECT 4.000 902.040 974.890 910.840 ;
        RECT 4.000 900.640 970.600 902.040 ;
        RECT 974.400 900.640 974.890 902.040 ;
        RECT 4.000 891.840 974.890 900.640 ;
        RECT 4.400 890.440 974.890 891.840 ;
        RECT 4.000 881.640 974.890 890.440 ;
        RECT 4.000 880.240 970.600 881.640 ;
        RECT 974.400 880.240 974.890 881.640 ;
        RECT 4.000 871.440 974.890 880.240 ;
        RECT 4.400 870.040 974.890 871.440 ;
        RECT 4.000 857.840 974.890 870.040 ;
        RECT 4.000 856.440 970.600 857.840 ;
        RECT 974.400 856.440 974.890 857.840 ;
        RECT 4.000 847.640 974.890 856.440 ;
        RECT 4.400 846.240 974.890 847.640 ;
        RECT 4.000 837.440 974.890 846.240 ;
        RECT 4.000 836.040 970.600 837.440 ;
        RECT 974.400 836.040 974.890 837.440 ;
        RECT 4.000 827.240 974.890 836.040 ;
        RECT 4.400 825.840 974.890 827.240 ;
        RECT 4.000 817.040 974.890 825.840 ;
        RECT 4.000 815.640 970.600 817.040 ;
        RECT 974.400 815.640 974.890 817.040 ;
        RECT 4.000 806.840 974.890 815.640 ;
        RECT 4.400 805.440 974.890 806.840 ;
        RECT 4.000 796.640 974.890 805.440 ;
        RECT 4.000 795.240 970.600 796.640 ;
        RECT 974.400 795.240 974.890 796.640 ;
        RECT 4.000 786.440 974.890 795.240 ;
        RECT 4.400 785.040 974.890 786.440 ;
        RECT 4.000 772.840 974.890 785.040 ;
        RECT 4.000 771.440 970.600 772.840 ;
        RECT 974.400 771.440 974.890 772.840 ;
        RECT 4.000 762.640 974.890 771.440 ;
        RECT 4.400 761.240 974.890 762.640 ;
        RECT 4.000 752.440 974.890 761.240 ;
        RECT 4.000 751.040 970.600 752.440 ;
        RECT 974.400 751.040 974.890 752.440 ;
        RECT 4.000 742.240 974.890 751.040 ;
        RECT 4.400 740.840 974.890 742.240 ;
        RECT 4.000 732.040 974.890 740.840 ;
        RECT 4.000 730.640 970.600 732.040 ;
        RECT 974.400 730.640 974.890 732.040 ;
        RECT 4.000 721.840 974.890 730.640 ;
        RECT 4.400 720.440 974.890 721.840 ;
        RECT 4.000 711.640 974.890 720.440 ;
        RECT 4.000 710.240 970.600 711.640 ;
        RECT 974.400 710.240 974.890 711.640 ;
        RECT 4.000 701.440 974.890 710.240 ;
        RECT 4.400 700.040 974.890 701.440 ;
        RECT 4.000 687.840 974.890 700.040 ;
        RECT 4.000 686.440 970.600 687.840 ;
        RECT 974.400 686.440 974.890 687.840 ;
        RECT 4.000 677.640 974.890 686.440 ;
        RECT 4.400 676.240 974.890 677.640 ;
        RECT 4.000 667.440 974.890 676.240 ;
        RECT 4.000 666.040 970.600 667.440 ;
        RECT 974.400 666.040 974.890 667.440 ;
        RECT 4.000 657.240 974.890 666.040 ;
        RECT 4.400 655.840 974.890 657.240 ;
        RECT 4.000 647.040 974.890 655.840 ;
        RECT 4.000 645.640 970.600 647.040 ;
        RECT 974.400 645.640 974.890 647.040 ;
        RECT 4.000 636.840 974.890 645.640 ;
        RECT 4.400 635.440 974.890 636.840 ;
        RECT 4.000 626.640 974.890 635.440 ;
        RECT 4.000 625.240 970.600 626.640 ;
        RECT 974.400 625.240 974.890 626.640 ;
        RECT 4.000 616.440 974.890 625.240 ;
        RECT 4.400 615.040 974.890 616.440 ;
        RECT 4.000 602.840 974.890 615.040 ;
        RECT 4.000 601.440 970.600 602.840 ;
        RECT 974.400 601.440 974.890 602.840 ;
        RECT 4.000 592.640 974.890 601.440 ;
        RECT 4.400 591.240 974.890 592.640 ;
        RECT 4.000 582.440 974.890 591.240 ;
        RECT 4.000 581.040 970.600 582.440 ;
        RECT 974.400 581.040 974.890 582.440 ;
        RECT 4.000 572.240 974.890 581.040 ;
        RECT 4.400 570.840 974.890 572.240 ;
        RECT 4.000 562.040 974.890 570.840 ;
        RECT 4.000 560.640 970.600 562.040 ;
        RECT 974.400 560.640 974.890 562.040 ;
        RECT 4.000 551.840 974.890 560.640 ;
        RECT 4.400 550.440 974.890 551.840 ;
        RECT 4.000 541.640 974.890 550.440 ;
        RECT 4.000 540.240 970.600 541.640 ;
        RECT 974.400 540.240 974.890 541.640 ;
        RECT 4.000 531.440 974.890 540.240 ;
        RECT 4.400 530.040 974.890 531.440 ;
        RECT 4.000 517.840 974.890 530.040 ;
        RECT 4.000 516.440 970.600 517.840 ;
        RECT 974.400 516.440 974.890 517.840 ;
        RECT 4.000 507.640 974.890 516.440 ;
        RECT 4.400 506.240 974.890 507.640 ;
        RECT 4.000 497.440 974.890 506.240 ;
        RECT 4.000 496.040 970.600 497.440 ;
        RECT 974.400 496.040 974.890 497.440 ;
        RECT 4.000 487.240 974.890 496.040 ;
        RECT 4.400 485.840 974.890 487.240 ;
        RECT 4.000 477.040 974.890 485.840 ;
        RECT 4.000 475.640 970.600 477.040 ;
        RECT 974.400 475.640 974.890 477.040 ;
        RECT 4.000 466.840 974.890 475.640 ;
        RECT 4.400 465.440 974.890 466.840 ;
        RECT 4.000 456.640 974.890 465.440 ;
        RECT 4.000 455.240 970.600 456.640 ;
        RECT 974.400 455.240 974.890 456.640 ;
        RECT 4.000 446.440 974.890 455.240 ;
        RECT 4.400 445.040 974.890 446.440 ;
        RECT 4.000 436.240 974.890 445.040 ;
        RECT 4.000 434.840 970.600 436.240 ;
        RECT 974.400 434.840 974.890 436.240 ;
        RECT 4.000 422.640 974.890 434.840 ;
        RECT 4.400 421.240 974.890 422.640 ;
        RECT 4.000 412.440 974.890 421.240 ;
        RECT 4.000 411.040 970.600 412.440 ;
        RECT 974.400 411.040 974.890 412.440 ;
        RECT 4.000 402.240 974.890 411.040 ;
        RECT 4.400 400.840 974.890 402.240 ;
        RECT 4.000 392.040 974.890 400.840 ;
        RECT 4.000 390.640 970.600 392.040 ;
        RECT 974.400 390.640 974.890 392.040 ;
        RECT 4.000 381.840 974.890 390.640 ;
        RECT 4.400 380.440 974.890 381.840 ;
        RECT 4.000 371.640 974.890 380.440 ;
        RECT 4.000 370.240 970.600 371.640 ;
        RECT 974.400 370.240 974.890 371.640 ;
        RECT 4.000 361.440 974.890 370.240 ;
        RECT 4.400 360.040 974.890 361.440 ;
        RECT 4.000 351.240 974.890 360.040 ;
        RECT 4.000 349.840 970.600 351.240 ;
        RECT 974.400 349.840 974.890 351.240 ;
        RECT 4.000 337.640 974.890 349.840 ;
        RECT 4.400 336.240 974.890 337.640 ;
        RECT 4.000 327.440 974.890 336.240 ;
        RECT 4.000 326.040 970.600 327.440 ;
        RECT 974.400 326.040 974.890 327.440 ;
        RECT 4.000 317.240 974.890 326.040 ;
        RECT 4.400 315.840 974.890 317.240 ;
        RECT 4.000 307.040 974.890 315.840 ;
        RECT 4.000 305.640 970.600 307.040 ;
        RECT 974.400 305.640 974.890 307.040 ;
        RECT 4.000 296.840 974.890 305.640 ;
        RECT 4.400 295.440 974.890 296.840 ;
        RECT 4.000 286.640 974.890 295.440 ;
        RECT 4.000 285.240 970.600 286.640 ;
        RECT 974.400 285.240 974.890 286.640 ;
        RECT 4.000 276.440 974.890 285.240 ;
        RECT 4.400 275.040 974.890 276.440 ;
        RECT 4.000 266.240 974.890 275.040 ;
        RECT 4.000 264.840 970.600 266.240 ;
        RECT 974.400 264.840 974.890 266.240 ;
        RECT 4.000 252.640 974.890 264.840 ;
        RECT 4.400 251.240 974.890 252.640 ;
        RECT 4.000 242.440 974.890 251.240 ;
        RECT 4.000 241.040 970.600 242.440 ;
        RECT 974.400 241.040 974.890 242.440 ;
        RECT 4.000 232.240 974.890 241.040 ;
        RECT 4.400 230.840 974.890 232.240 ;
        RECT 4.000 222.040 974.890 230.840 ;
        RECT 4.000 220.640 970.600 222.040 ;
        RECT 974.400 220.640 974.890 222.040 ;
        RECT 4.000 211.840 974.890 220.640 ;
        RECT 4.400 210.440 974.890 211.840 ;
        RECT 4.000 201.640 974.890 210.440 ;
        RECT 4.000 200.240 970.600 201.640 ;
        RECT 974.400 200.240 974.890 201.640 ;
        RECT 4.000 191.440 974.890 200.240 ;
        RECT 4.400 190.040 974.890 191.440 ;
        RECT 4.000 181.240 974.890 190.040 ;
        RECT 4.000 179.840 970.600 181.240 ;
        RECT 974.400 179.840 974.890 181.240 ;
        RECT 4.000 167.640 974.890 179.840 ;
        RECT 4.400 166.240 974.890 167.640 ;
        RECT 4.000 157.440 974.890 166.240 ;
        RECT 4.000 156.040 970.600 157.440 ;
        RECT 974.400 156.040 974.890 157.440 ;
        RECT 4.000 147.240 974.890 156.040 ;
        RECT 4.400 145.840 974.890 147.240 ;
        RECT 4.000 137.040 974.890 145.840 ;
        RECT 4.000 135.640 970.600 137.040 ;
        RECT 974.400 135.640 974.890 137.040 ;
        RECT 4.000 126.840 974.890 135.640 ;
        RECT 4.400 125.440 974.890 126.840 ;
        RECT 4.000 116.640 974.890 125.440 ;
        RECT 4.000 115.240 970.600 116.640 ;
        RECT 974.400 115.240 974.890 116.640 ;
        RECT 4.000 106.440 974.890 115.240 ;
        RECT 4.400 105.040 974.890 106.440 ;
        RECT 4.000 96.240 974.890 105.040 ;
        RECT 4.000 94.840 970.600 96.240 ;
        RECT 974.400 94.840 974.890 96.240 ;
        RECT 4.000 82.640 974.890 94.840 ;
        RECT 4.400 81.240 974.890 82.640 ;
        RECT 4.000 72.440 974.890 81.240 ;
        RECT 4.000 71.040 970.600 72.440 ;
        RECT 974.400 71.040 974.890 72.440 ;
        RECT 4.000 62.240 974.890 71.040 ;
        RECT 4.400 60.840 974.890 62.240 ;
        RECT 4.000 52.040 974.890 60.840 ;
        RECT 4.000 50.640 970.600 52.040 ;
        RECT 974.400 50.640 974.890 52.040 ;
        RECT 4.000 41.840 974.890 50.640 ;
        RECT 4.400 40.440 974.890 41.840 ;
        RECT 4.000 31.640 974.890 40.440 ;
        RECT 4.000 30.240 970.600 31.640 ;
        RECT 974.400 30.240 974.890 31.640 ;
        RECT 4.000 21.440 974.890 30.240 ;
        RECT 4.400 20.040 974.890 21.440 ;
        RECT 4.000 11.240 974.890 20.040 ;
        RECT 4.000 10.390 970.600 11.240 ;
        RECT 974.400 10.390 974.890 11.240 ;
      LAYER met4 ;
        RECT 85.855 11.735 97.440 1886.825 ;
        RECT 99.840 11.735 174.240 1886.825 ;
        RECT 176.640 11.735 251.040 1886.825 ;
        RECT 253.440 11.735 327.840 1886.825 ;
        RECT 330.240 11.735 404.640 1886.825 ;
        RECT 407.040 11.735 481.440 1886.825 ;
        RECT 483.840 11.735 558.240 1886.825 ;
        RECT 560.640 11.735 635.040 1886.825 ;
        RECT 637.440 11.735 711.840 1886.825 ;
        RECT 714.240 11.735 788.640 1886.825 ;
        RECT 791.040 11.735 865.440 1886.825 ;
        RECT 867.840 11.735 906.825 1886.825 ;
  END
END Top_Module_4_ALU
END LIBRARY

