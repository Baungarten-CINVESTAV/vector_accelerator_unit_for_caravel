magic
tech sky130A
magscale 1 2
timestamp 1676901211
<< obsli1 >>
rect 1104 2159 193844 377553
<< obsm1 >>
rect 14 2128 194934 377584
<< metal2 >>
rect 1950 379200 2006 379800
rect 5814 379200 5870 379800
rect 9678 379200 9734 379800
rect 13542 379200 13598 379800
rect 18050 379200 18106 379800
rect 21914 379200 21970 379800
rect 25778 379200 25834 379800
rect 29642 379200 29698 379800
rect 34150 379200 34206 379800
rect 38014 379200 38070 379800
rect 41878 379200 41934 379800
rect 45742 379200 45798 379800
rect 50250 379200 50306 379800
rect 54114 379200 54170 379800
rect 57978 379200 58034 379800
rect 61842 379200 61898 379800
rect 66350 379200 66406 379800
rect 70214 379200 70270 379800
rect 74078 379200 74134 379800
rect 77942 379200 77998 379800
rect 82450 379200 82506 379800
rect 86314 379200 86370 379800
rect 90178 379200 90234 379800
rect 94042 379200 94098 379800
rect 98550 379200 98606 379800
rect 102414 379200 102470 379800
rect 106278 379200 106334 379800
rect 110142 379200 110198 379800
rect 114650 379200 114706 379800
rect 118514 379200 118570 379800
rect 122378 379200 122434 379800
rect 126242 379200 126298 379800
rect 130750 379200 130806 379800
rect 134614 379200 134670 379800
rect 138478 379200 138534 379800
rect 142342 379200 142398 379800
rect 146850 379200 146906 379800
rect 150714 379200 150770 379800
rect 154578 379200 154634 379800
rect 158442 379200 158498 379800
rect 162950 379200 163006 379800
rect 166814 379200 166870 379800
rect 170678 379200 170734 379800
rect 174542 379200 174598 379800
rect 179050 379200 179106 379800
rect 182914 379200 182970 379800
rect 186778 379200 186834 379800
rect 190642 379200 190698 379800
rect 194506 379200 194562 379800
rect 18 200 74 800
rect 3882 200 3938 800
rect 7746 200 7802 800
rect 11610 200 11666 800
rect 15474 200 15530 800
rect 19982 200 20038 800
rect 23846 200 23902 800
rect 27710 200 27766 800
rect 31574 200 31630 800
rect 36082 200 36138 800
rect 39946 200 40002 800
rect 43810 200 43866 800
rect 47674 200 47730 800
rect 52182 200 52238 800
rect 56046 200 56102 800
rect 59910 200 59966 800
rect 63774 200 63830 800
rect 68282 200 68338 800
rect 72146 200 72202 800
rect 76010 200 76066 800
rect 79874 200 79930 800
rect 84382 200 84438 800
rect 88246 200 88302 800
rect 92110 200 92166 800
rect 95974 200 96030 800
rect 100482 200 100538 800
rect 104346 200 104402 800
rect 108210 200 108266 800
rect 112074 200 112130 800
rect 116582 200 116638 800
rect 120446 200 120502 800
rect 124310 200 124366 800
rect 128174 200 128230 800
rect 132682 200 132738 800
rect 136546 200 136602 800
rect 140410 200 140466 800
rect 144274 200 144330 800
rect 148782 200 148838 800
rect 152646 200 152702 800
rect 156510 200 156566 800
rect 160374 200 160430 800
rect 164882 200 164938 800
rect 168746 200 168802 800
rect 172610 200 172666 800
rect 176474 200 176530 800
rect 180982 200 181038 800
rect 184846 200 184902 800
rect 188710 200 188766 800
rect 192574 200 192630 800
<< obsm2 >>
rect 20 379144 1894 379200
rect 2062 379144 5758 379200
rect 5926 379144 9622 379200
rect 9790 379144 13486 379200
rect 13654 379144 17994 379200
rect 18162 379144 21858 379200
rect 22026 379144 25722 379200
rect 25890 379144 29586 379200
rect 29754 379144 34094 379200
rect 34262 379144 37958 379200
rect 38126 379144 41822 379200
rect 41990 379144 45686 379200
rect 45854 379144 50194 379200
rect 50362 379144 54058 379200
rect 54226 379144 57922 379200
rect 58090 379144 61786 379200
rect 61954 379144 66294 379200
rect 66462 379144 70158 379200
rect 70326 379144 74022 379200
rect 74190 379144 77886 379200
rect 78054 379144 82394 379200
rect 82562 379144 86258 379200
rect 86426 379144 90122 379200
rect 90290 379144 93986 379200
rect 94154 379144 98494 379200
rect 98662 379144 102358 379200
rect 102526 379144 106222 379200
rect 106390 379144 110086 379200
rect 110254 379144 114594 379200
rect 114762 379144 118458 379200
rect 118626 379144 122322 379200
rect 122490 379144 126186 379200
rect 126354 379144 130694 379200
rect 130862 379144 134558 379200
rect 134726 379144 138422 379200
rect 138590 379144 142286 379200
rect 142454 379144 146794 379200
rect 146962 379144 150658 379200
rect 150826 379144 154522 379200
rect 154690 379144 158386 379200
rect 158554 379144 162894 379200
rect 163062 379144 166758 379200
rect 166926 379144 170622 379200
rect 170790 379144 174486 379200
rect 174654 379144 178994 379200
rect 179162 379144 182858 379200
rect 183026 379144 186722 379200
rect 186890 379144 190586 379200
rect 190754 379144 194450 379200
rect 194618 379144 194930 379200
rect 20 856 194930 379144
rect 130 734 3826 856
rect 3994 734 7690 856
rect 7858 734 11554 856
rect 11722 734 15418 856
rect 15586 734 19926 856
rect 20094 734 23790 856
rect 23958 734 27654 856
rect 27822 734 31518 856
rect 31686 734 36026 856
rect 36194 734 39890 856
rect 40058 734 43754 856
rect 43922 734 47618 856
rect 47786 734 52126 856
rect 52294 734 55990 856
rect 56158 734 59854 856
rect 60022 734 63718 856
rect 63886 734 68226 856
rect 68394 734 72090 856
rect 72258 734 75954 856
rect 76122 734 79818 856
rect 79986 734 84326 856
rect 84494 734 88190 856
rect 88358 734 92054 856
rect 92222 734 95918 856
rect 96086 734 100426 856
rect 100594 734 104290 856
rect 104458 734 108154 856
rect 108322 734 112018 856
rect 112186 734 116526 856
rect 116694 734 120390 856
rect 120558 734 124254 856
rect 124422 734 128118 856
rect 128286 734 132626 856
rect 132794 734 136490 856
rect 136658 734 140354 856
rect 140522 734 144218 856
rect 144386 734 148726 856
rect 148894 734 152590 856
rect 152758 734 156454 856
rect 156622 734 160318 856
rect 160486 734 164826 856
rect 164994 734 168690 856
rect 168858 734 172554 856
rect 172722 734 176418 856
rect 176586 734 180926 856
rect 181094 734 184790 856
rect 184958 734 188654 856
rect 188822 734 192518 856
rect 192686 734 194930 856
<< metal3 >>
rect 200 377408 800 377528
rect 194200 375368 194800 375488
rect 200 373328 800 373448
rect 194200 371288 194800 371408
rect 200 369248 800 369368
rect 194200 367208 194800 367328
rect 200 365168 800 365288
rect 194200 363128 194800 363248
rect 200 360408 800 360528
rect 194200 358368 194800 358488
rect 200 356328 800 356448
rect 194200 354288 194800 354408
rect 200 352248 800 352368
rect 194200 350208 194800 350328
rect 200 348168 800 348288
rect 194200 346128 194800 346248
rect 200 343408 800 343528
rect 194200 341368 194800 341488
rect 200 339328 800 339448
rect 194200 337288 194800 337408
rect 200 335248 800 335368
rect 194200 333208 194800 333328
rect 200 331168 800 331288
rect 194200 329128 194800 329248
rect 200 326408 800 326528
rect 194200 324368 194800 324488
rect 200 322328 800 322448
rect 194200 320288 194800 320408
rect 200 318248 800 318368
rect 194200 316208 194800 316328
rect 200 314168 800 314288
rect 194200 312128 194800 312248
rect 200 309408 800 309528
rect 194200 307368 194800 307488
rect 200 305328 800 305448
rect 194200 303288 194800 303408
rect 200 301248 800 301368
rect 194200 299208 194800 299328
rect 200 297168 800 297288
rect 194200 295128 194800 295248
rect 200 292408 800 292528
rect 194200 290368 194800 290488
rect 200 288328 800 288448
rect 194200 286288 194800 286408
rect 200 284248 800 284368
rect 194200 282208 194800 282328
rect 200 280168 800 280288
rect 194200 278128 194800 278248
rect 200 276088 800 276208
rect 194200 273368 194800 273488
rect 200 271328 800 271448
rect 194200 269288 194800 269408
rect 200 267248 800 267368
rect 194200 265208 194800 265328
rect 200 263168 800 263288
rect 194200 261128 194800 261248
rect 200 259088 800 259208
rect 194200 256368 194800 256488
rect 200 254328 800 254448
rect 194200 252288 194800 252408
rect 200 250248 800 250368
rect 194200 248208 194800 248328
rect 200 246168 800 246288
rect 194200 244128 194800 244248
rect 200 242088 800 242208
rect 194200 239368 194800 239488
rect 200 237328 800 237448
rect 194200 235288 194800 235408
rect 200 233248 800 233368
rect 194200 231208 194800 231328
rect 200 229168 800 229288
rect 194200 227128 194800 227248
rect 200 225088 800 225208
rect 194200 222368 194800 222488
rect 200 220328 800 220448
rect 194200 218288 194800 218408
rect 200 216248 800 216368
rect 194200 214208 194800 214328
rect 200 212168 800 212288
rect 194200 210128 194800 210248
rect 200 208088 800 208208
rect 194200 205368 194800 205488
rect 200 203328 800 203448
rect 194200 201288 194800 201408
rect 200 199248 800 199368
rect 194200 197208 194800 197328
rect 200 195168 800 195288
rect 194200 193128 194800 193248
rect 200 191088 800 191208
rect 194200 188368 194800 188488
rect 200 186328 800 186448
rect 194200 184288 194800 184408
rect 200 182248 800 182368
rect 194200 180208 194800 180328
rect 200 178168 800 178288
rect 194200 176128 194800 176248
rect 200 174088 800 174208
rect 194200 171368 194800 171488
rect 200 169328 800 169448
rect 194200 167288 194800 167408
rect 200 165248 800 165368
rect 194200 163208 194800 163328
rect 200 161168 800 161288
rect 194200 159128 194800 159248
rect 200 157088 800 157208
rect 194200 154368 194800 154488
rect 200 152328 800 152448
rect 194200 150288 194800 150408
rect 200 148248 800 148368
rect 194200 146208 194800 146328
rect 200 144168 800 144288
rect 194200 142128 194800 142248
rect 200 140088 800 140208
rect 194200 137368 194800 137488
rect 200 135328 800 135448
rect 194200 133288 194800 133408
rect 200 131248 800 131368
rect 194200 129208 194800 129328
rect 200 127168 800 127288
rect 194200 125128 194800 125248
rect 200 123088 800 123208
rect 194200 120368 194800 120488
rect 200 118328 800 118448
rect 194200 116288 194800 116408
rect 200 114248 800 114368
rect 194200 112208 194800 112328
rect 200 110168 800 110288
rect 194200 108128 194800 108248
rect 200 106088 800 106208
rect 194200 103368 194800 103488
rect 200 101328 800 101448
rect 194200 99288 194800 99408
rect 200 97248 800 97368
rect 194200 95208 194800 95328
rect 200 93168 800 93288
rect 194200 91128 194800 91248
rect 200 89088 800 89208
rect 194200 87048 194800 87168
rect 200 84328 800 84448
rect 194200 82288 194800 82408
rect 200 80248 800 80368
rect 194200 78208 194800 78328
rect 200 76168 800 76288
rect 194200 74128 194800 74248
rect 200 72088 800 72208
rect 194200 70048 194800 70168
rect 200 67328 800 67448
rect 194200 65288 194800 65408
rect 200 63248 800 63368
rect 194200 61208 194800 61328
rect 200 59168 800 59288
rect 194200 57128 194800 57248
rect 200 55088 800 55208
rect 194200 53048 194800 53168
rect 200 50328 800 50448
rect 194200 48288 194800 48408
rect 200 46248 800 46368
rect 194200 44208 194800 44328
rect 200 42168 800 42288
rect 194200 40128 194800 40248
rect 200 38088 800 38208
rect 194200 36048 194800 36168
rect 200 33328 800 33448
rect 194200 31288 194800 31408
rect 200 29248 800 29368
rect 194200 27208 194800 27328
rect 200 25168 800 25288
rect 194200 23128 194800 23248
rect 200 21088 800 21208
rect 194200 19048 194800 19168
rect 200 16328 800 16448
rect 194200 14288 194800 14408
rect 200 12248 800 12368
rect 194200 10208 194800 10328
rect 200 8168 800 8288
rect 194200 6128 194800 6248
rect 200 4088 800 4208
rect 194200 2048 194800 2168
<< obsm3 >>
rect 880 377328 194978 377569
rect 800 375568 194978 377328
rect 800 375288 194120 375568
rect 194880 375288 194978 375568
rect 800 373528 194978 375288
rect 880 373248 194978 373528
rect 800 371488 194978 373248
rect 800 371208 194120 371488
rect 194880 371208 194978 371488
rect 800 369448 194978 371208
rect 880 369168 194978 369448
rect 800 367408 194978 369168
rect 800 367128 194120 367408
rect 194880 367128 194978 367408
rect 800 365368 194978 367128
rect 880 365088 194978 365368
rect 800 363328 194978 365088
rect 800 363048 194120 363328
rect 194880 363048 194978 363328
rect 800 360608 194978 363048
rect 880 360328 194978 360608
rect 800 358568 194978 360328
rect 800 358288 194120 358568
rect 194880 358288 194978 358568
rect 800 356528 194978 358288
rect 880 356248 194978 356528
rect 800 354488 194978 356248
rect 800 354208 194120 354488
rect 194880 354208 194978 354488
rect 800 352448 194978 354208
rect 880 352168 194978 352448
rect 800 350408 194978 352168
rect 800 350128 194120 350408
rect 194880 350128 194978 350408
rect 800 348368 194978 350128
rect 880 348088 194978 348368
rect 800 346328 194978 348088
rect 800 346048 194120 346328
rect 194880 346048 194978 346328
rect 800 343608 194978 346048
rect 880 343328 194978 343608
rect 800 341568 194978 343328
rect 800 341288 194120 341568
rect 194880 341288 194978 341568
rect 800 339528 194978 341288
rect 880 339248 194978 339528
rect 800 337488 194978 339248
rect 800 337208 194120 337488
rect 194880 337208 194978 337488
rect 800 335448 194978 337208
rect 880 335168 194978 335448
rect 800 333408 194978 335168
rect 800 333128 194120 333408
rect 194880 333128 194978 333408
rect 800 331368 194978 333128
rect 880 331088 194978 331368
rect 800 329328 194978 331088
rect 800 329048 194120 329328
rect 194880 329048 194978 329328
rect 800 326608 194978 329048
rect 880 326328 194978 326608
rect 800 324568 194978 326328
rect 800 324288 194120 324568
rect 194880 324288 194978 324568
rect 800 322528 194978 324288
rect 880 322248 194978 322528
rect 800 320488 194978 322248
rect 800 320208 194120 320488
rect 194880 320208 194978 320488
rect 800 318448 194978 320208
rect 880 318168 194978 318448
rect 800 316408 194978 318168
rect 800 316128 194120 316408
rect 194880 316128 194978 316408
rect 800 314368 194978 316128
rect 880 314088 194978 314368
rect 800 312328 194978 314088
rect 800 312048 194120 312328
rect 194880 312048 194978 312328
rect 800 309608 194978 312048
rect 880 309328 194978 309608
rect 800 307568 194978 309328
rect 800 307288 194120 307568
rect 194880 307288 194978 307568
rect 800 305528 194978 307288
rect 880 305248 194978 305528
rect 800 303488 194978 305248
rect 800 303208 194120 303488
rect 194880 303208 194978 303488
rect 800 301448 194978 303208
rect 880 301168 194978 301448
rect 800 299408 194978 301168
rect 800 299128 194120 299408
rect 194880 299128 194978 299408
rect 800 297368 194978 299128
rect 880 297088 194978 297368
rect 800 295328 194978 297088
rect 800 295048 194120 295328
rect 194880 295048 194978 295328
rect 800 292608 194978 295048
rect 880 292328 194978 292608
rect 800 290568 194978 292328
rect 800 290288 194120 290568
rect 194880 290288 194978 290568
rect 800 288528 194978 290288
rect 880 288248 194978 288528
rect 800 286488 194978 288248
rect 800 286208 194120 286488
rect 194880 286208 194978 286488
rect 800 284448 194978 286208
rect 880 284168 194978 284448
rect 800 282408 194978 284168
rect 800 282128 194120 282408
rect 194880 282128 194978 282408
rect 800 280368 194978 282128
rect 880 280088 194978 280368
rect 800 278328 194978 280088
rect 800 278048 194120 278328
rect 194880 278048 194978 278328
rect 800 276288 194978 278048
rect 880 276008 194978 276288
rect 800 273568 194978 276008
rect 800 273288 194120 273568
rect 194880 273288 194978 273568
rect 800 271528 194978 273288
rect 880 271248 194978 271528
rect 800 269488 194978 271248
rect 800 269208 194120 269488
rect 194880 269208 194978 269488
rect 800 267448 194978 269208
rect 880 267168 194978 267448
rect 800 265408 194978 267168
rect 800 265128 194120 265408
rect 194880 265128 194978 265408
rect 800 263368 194978 265128
rect 880 263088 194978 263368
rect 800 261328 194978 263088
rect 800 261048 194120 261328
rect 194880 261048 194978 261328
rect 800 259288 194978 261048
rect 880 259008 194978 259288
rect 800 256568 194978 259008
rect 800 256288 194120 256568
rect 194880 256288 194978 256568
rect 800 254528 194978 256288
rect 880 254248 194978 254528
rect 800 252488 194978 254248
rect 800 252208 194120 252488
rect 194880 252208 194978 252488
rect 800 250448 194978 252208
rect 880 250168 194978 250448
rect 800 248408 194978 250168
rect 800 248128 194120 248408
rect 194880 248128 194978 248408
rect 800 246368 194978 248128
rect 880 246088 194978 246368
rect 800 244328 194978 246088
rect 800 244048 194120 244328
rect 194880 244048 194978 244328
rect 800 242288 194978 244048
rect 880 242008 194978 242288
rect 800 239568 194978 242008
rect 800 239288 194120 239568
rect 194880 239288 194978 239568
rect 800 237528 194978 239288
rect 880 237248 194978 237528
rect 800 235488 194978 237248
rect 800 235208 194120 235488
rect 194880 235208 194978 235488
rect 800 233448 194978 235208
rect 880 233168 194978 233448
rect 800 231408 194978 233168
rect 800 231128 194120 231408
rect 194880 231128 194978 231408
rect 800 229368 194978 231128
rect 880 229088 194978 229368
rect 800 227328 194978 229088
rect 800 227048 194120 227328
rect 194880 227048 194978 227328
rect 800 225288 194978 227048
rect 880 225008 194978 225288
rect 800 222568 194978 225008
rect 800 222288 194120 222568
rect 194880 222288 194978 222568
rect 800 220528 194978 222288
rect 880 220248 194978 220528
rect 800 218488 194978 220248
rect 800 218208 194120 218488
rect 194880 218208 194978 218488
rect 800 216448 194978 218208
rect 880 216168 194978 216448
rect 800 214408 194978 216168
rect 800 214128 194120 214408
rect 194880 214128 194978 214408
rect 800 212368 194978 214128
rect 880 212088 194978 212368
rect 800 210328 194978 212088
rect 800 210048 194120 210328
rect 194880 210048 194978 210328
rect 800 208288 194978 210048
rect 880 208008 194978 208288
rect 800 205568 194978 208008
rect 800 205288 194120 205568
rect 194880 205288 194978 205568
rect 800 203528 194978 205288
rect 880 203248 194978 203528
rect 800 201488 194978 203248
rect 800 201208 194120 201488
rect 194880 201208 194978 201488
rect 800 199448 194978 201208
rect 880 199168 194978 199448
rect 800 197408 194978 199168
rect 800 197128 194120 197408
rect 194880 197128 194978 197408
rect 800 195368 194978 197128
rect 880 195088 194978 195368
rect 800 193328 194978 195088
rect 800 193048 194120 193328
rect 194880 193048 194978 193328
rect 800 191288 194978 193048
rect 880 191008 194978 191288
rect 800 188568 194978 191008
rect 800 188288 194120 188568
rect 194880 188288 194978 188568
rect 800 186528 194978 188288
rect 880 186248 194978 186528
rect 800 184488 194978 186248
rect 800 184208 194120 184488
rect 194880 184208 194978 184488
rect 800 182448 194978 184208
rect 880 182168 194978 182448
rect 800 180408 194978 182168
rect 800 180128 194120 180408
rect 194880 180128 194978 180408
rect 800 178368 194978 180128
rect 880 178088 194978 178368
rect 800 176328 194978 178088
rect 800 176048 194120 176328
rect 194880 176048 194978 176328
rect 800 174288 194978 176048
rect 880 174008 194978 174288
rect 800 171568 194978 174008
rect 800 171288 194120 171568
rect 194880 171288 194978 171568
rect 800 169528 194978 171288
rect 880 169248 194978 169528
rect 800 167488 194978 169248
rect 800 167208 194120 167488
rect 194880 167208 194978 167488
rect 800 165448 194978 167208
rect 880 165168 194978 165448
rect 800 163408 194978 165168
rect 800 163128 194120 163408
rect 194880 163128 194978 163408
rect 800 161368 194978 163128
rect 880 161088 194978 161368
rect 800 159328 194978 161088
rect 800 159048 194120 159328
rect 194880 159048 194978 159328
rect 800 157288 194978 159048
rect 880 157008 194978 157288
rect 800 154568 194978 157008
rect 800 154288 194120 154568
rect 194880 154288 194978 154568
rect 800 152528 194978 154288
rect 880 152248 194978 152528
rect 800 150488 194978 152248
rect 800 150208 194120 150488
rect 194880 150208 194978 150488
rect 800 148448 194978 150208
rect 880 148168 194978 148448
rect 800 146408 194978 148168
rect 800 146128 194120 146408
rect 194880 146128 194978 146408
rect 800 144368 194978 146128
rect 880 144088 194978 144368
rect 800 142328 194978 144088
rect 800 142048 194120 142328
rect 194880 142048 194978 142328
rect 800 140288 194978 142048
rect 880 140008 194978 140288
rect 800 137568 194978 140008
rect 800 137288 194120 137568
rect 194880 137288 194978 137568
rect 800 135528 194978 137288
rect 880 135248 194978 135528
rect 800 133488 194978 135248
rect 800 133208 194120 133488
rect 194880 133208 194978 133488
rect 800 131448 194978 133208
rect 880 131168 194978 131448
rect 800 129408 194978 131168
rect 800 129128 194120 129408
rect 194880 129128 194978 129408
rect 800 127368 194978 129128
rect 880 127088 194978 127368
rect 800 125328 194978 127088
rect 800 125048 194120 125328
rect 194880 125048 194978 125328
rect 800 123288 194978 125048
rect 880 123008 194978 123288
rect 800 120568 194978 123008
rect 800 120288 194120 120568
rect 194880 120288 194978 120568
rect 800 118528 194978 120288
rect 880 118248 194978 118528
rect 800 116488 194978 118248
rect 800 116208 194120 116488
rect 194880 116208 194978 116488
rect 800 114448 194978 116208
rect 880 114168 194978 114448
rect 800 112408 194978 114168
rect 800 112128 194120 112408
rect 194880 112128 194978 112408
rect 800 110368 194978 112128
rect 880 110088 194978 110368
rect 800 108328 194978 110088
rect 800 108048 194120 108328
rect 194880 108048 194978 108328
rect 800 106288 194978 108048
rect 880 106008 194978 106288
rect 800 103568 194978 106008
rect 800 103288 194120 103568
rect 194880 103288 194978 103568
rect 800 101528 194978 103288
rect 880 101248 194978 101528
rect 800 99488 194978 101248
rect 800 99208 194120 99488
rect 194880 99208 194978 99488
rect 800 97448 194978 99208
rect 880 97168 194978 97448
rect 800 95408 194978 97168
rect 800 95128 194120 95408
rect 194880 95128 194978 95408
rect 800 93368 194978 95128
rect 880 93088 194978 93368
rect 800 91328 194978 93088
rect 800 91048 194120 91328
rect 194880 91048 194978 91328
rect 800 89288 194978 91048
rect 880 89008 194978 89288
rect 800 87248 194978 89008
rect 800 86968 194120 87248
rect 194880 86968 194978 87248
rect 800 84528 194978 86968
rect 880 84248 194978 84528
rect 800 82488 194978 84248
rect 800 82208 194120 82488
rect 194880 82208 194978 82488
rect 800 80448 194978 82208
rect 880 80168 194978 80448
rect 800 78408 194978 80168
rect 800 78128 194120 78408
rect 194880 78128 194978 78408
rect 800 76368 194978 78128
rect 880 76088 194978 76368
rect 800 74328 194978 76088
rect 800 74048 194120 74328
rect 194880 74048 194978 74328
rect 800 72288 194978 74048
rect 880 72008 194978 72288
rect 800 70248 194978 72008
rect 800 69968 194120 70248
rect 194880 69968 194978 70248
rect 800 67528 194978 69968
rect 880 67248 194978 67528
rect 800 65488 194978 67248
rect 800 65208 194120 65488
rect 194880 65208 194978 65488
rect 800 63448 194978 65208
rect 880 63168 194978 63448
rect 800 61408 194978 63168
rect 800 61128 194120 61408
rect 194880 61128 194978 61408
rect 800 59368 194978 61128
rect 880 59088 194978 59368
rect 800 57328 194978 59088
rect 800 57048 194120 57328
rect 194880 57048 194978 57328
rect 800 55288 194978 57048
rect 880 55008 194978 55288
rect 800 53248 194978 55008
rect 800 52968 194120 53248
rect 194880 52968 194978 53248
rect 800 50528 194978 52968
rect 880 50248 194978 50528
rect 800 48488 194978 50248
rect 800 48208 194120 48488
rect 194880 48208 194978 48488
rect 800 46448 194978 48208
rect 880 46168 194978 46448
rect 800 44408 194978 46168
rect 800 44128 194120 44408
rect 194880 44128 194978 44408
rect 800 42368 194978 44128
rect 880 42088 194978 42368
rect 800 40328 194978 42088
rect 800 40048 194120 40328
rect 194880 40048 194978 40328
rect 800 38288 194978 40048
rect 880 38008 194978 38288
rect 800 36248 194978 38008
rect 800 35968 194120 36248
rect 194880 35968 194978 36248
rect 800 33528 194978 35968
rect 880 33248 194978 33528
rect 800 31488 194978 33248
rect 800 31208 194120 31488
rect 194880 31208 194978 31488
rect 800 29448 194978 31208
rect 880 29168 194978 29448
rect 800 27408 194978 29168
rect 800 27128 194120 27408
rect 194880 27128 194978 27408
rect 800 25368 194978 27128
rect 880 25088 194978 25368
rect 800 23328 194978 25088
rect 800 23048 194120 23328
rect 194880 23048 194978 23328
rect 800 21288 194978 23048
rect 880 21008 194978 21288
rect 800 19248 194978 21008
rect 800 18968 194120 19248
rect 194880 18968 194978 19248
rect 800 16528 194978 18968
rect 880 16248 194978 16528
rect 800 14488 194978 16248
rect 800 14208 194120 14488
rect 194880 14208 194978 14488
rect 800 12448 194978 14208
rect 880 12168 194978 12448
rect 800 10408 194978 12168
rect 800 10128 194120 10408
rect 194880 10128 194978 10408
rect 800 8368 194978 10128
rect 880 8088 194978 8368
rect 800 6328 194978 8088
rect 800 6048 194120 6328
rect 194880 6048 194978 6328
rect 800 4288 194978 6048
rect 880 4008 194978 4288
rect 800 2248 194978 4008
rect 800 2078 194120 2248
rect 194880 2078 194978 2248
<< metal4 >>
rect 4208 2128 4528 377584
rect 19568 2128 19888 377584
rect 34928 2128 35248 377584
rect 50288 2128 50608 377584
rect 65648 2128 65968 377584
rect 81008 2128 81328 377584
rect 96368 2128 96688 377584
rect 111728 2128 112048 377584
rect 127088 2128 127408 377584
rect 142448 2128 142768 377584
rect 157808 2128 158128 377584
rect 173168 2128 173488 377584
rect 188528 2128 188848 377584
<< obsm4 >>
rect 17171 2347 19488 377365
rect 19968 2347 34848 377365
rect 35328 2347 50208 377365
rect 50688 2347 65568 377365
rect 66048 2347 80928 377365
rect 81408 2347 96288 377365
rect 96768 2347 111648 377365
rect 112128 2347 127008 377365
rect 127488 2347 142368 377365
rect 142848 2347 157728 377365
rect 158208 2347 173088 377365
rect 173568 2347 181365 377365
<< labels >>
rlabel metal2 s 186778 379200 186834 379800 6 ALU_Output[0]
port 1 nsew signal output
rlabel metal3 s 200 267248 800 267368 6 ALU_Output[100]
port 2 nsew signal output
rlabel metal3 s 194200 23128 194800 23248 6 ALU_Output[101]
port 3 nsew signal output
rlabel metal3 s 194200 341368 194800 341488 6 ALU_Output[102]
port 4 nsew signal output
rlabel metal2 s 41878 379200 41934 379800 6 ALU_Output[103]
port 5 nsew signal output
rlabel metal3 s 194200 116288 194800 116408 6 ALU_Output[104]
port 6 nsew signal output
rlabel metal3 s 194200 337288 194800 337408 6 ALU_Output[105]
port 7 nsew signal output
rlabel metal2 s 118514 379200 118570 379800 6 ALU_Output[106]
port 8 nsew signal output
rlabel metal3 s 200 263168 800 263288 6 ALU_Output[107]
port 9 nsew signal output
rlabel metal3 s 194200 44208 194800 44328 6 ALU_Output[108]
port 10 nsew signal output
rlabel metal3 s 200 208088 800 208208 6 ALU_Output[109]
port 11 nsew signal output
rlabel metal3 s 200 8168 800 8288 6 ALU_Output[10]
port 12 nsew signal output
rlabel metal2 s 114650 379200 114706 379800 6 ALU_Output[110]
port 13 nsew signal output
rlabel metal3 s 194200 214208 194800 214328 6 ALU_Output[111]
port 14 nsew signal output
rlabel metal3 s 200 297168 800 297288 6 ALU_Output[112]
port 15 nsew signal output
rlabel metal3 s 200 352248 800 352368 6 ALU_Output[113]
port 16 nsew signal output
rlabel metal3 s 194200 61208 194800 61328 6 ALU_Output[114]
port 17 nsew signal output
rlabel metal3 s 200 229168 800 229288 6 ALU_Output[115]
port 18 nsew signal output
rlabel metal3 s 194200 65288 194800 65408 6 ALU_Output[116]
port 19 nsew signal output
rlabel metal2 s 95974 200 96030 800 6 ALU_Output[117]
port 20 nsew signal output
rlabel metal2 s 130750 379200 130806 379800 6 ALU_Output[118]
port 21 nsew signal output
rlabel metal2 s 72146 200 72202 800 6 ALU_Output[119]
port 22 nsew signal output
rlabel metal2 s 54114 379200 54170 379800 6 ALU_Output[11]
port 23 nsew signal output
rlabel metal3 s 200 318248 800 318368 6 ALU_Output[120]
port 24 nsew signal output
rlabel metal3 s 200 259088 800 259208 6 ALU_Output[121]
port 25 nsew signal output
rlabel metal3 s 200 216248 800 216368 6 ALU_Output[122]
port 26 nsew signal output
rlabel metal3 s 200 97248 800 97368 6 ALU_Output[123]
port 27 nsew signal output
rlabel metal3 s 194200 256368 194800 256488 6 ALU_Output[124]
port 28 nsew signal output
rlabel metal2 s 50250 379200 50306 379800 6 ALU_Output[125]
port 29 nsew signal output
rlabel metal3 s 200 199248 800 199368 6 ALU_Output[126]
port 30 nsew signal output
rlabel metal2 s 112074 200 112130 800 6 ALU_Output[127]
port 31 nsew signal output
rlabel metal3 s 194200 261128 194800 261248 6 ALU_Output[12]
port 32 nsew signal output
rlabel metal2 s 5814 379200 5870 379800 6 ALU_Output[13]
port 33 nsew signal output
rlabel metal3 s 194200 82288 194800 82408 6 ALU_Output[14]
port 34 nsew signal output
rlabel metal3 s 194200 14288 194800 14408 6 ALU_Output[15]
port 35 nsew signal output
rlabel metal2 s 116582 200 116638 800 6 ALU_Output[16]
port 36 nsew signal output
rlabel metal3 s 200 246168 800 246288 6 ALU_Output[17]
port 37 nsew signal output
rlabel metal3 s 200 225088 800 225208 6 ALU_Output[18]
port 38 nsew signal output
rlabel metal3 s 194200 31288 194800 31408 6 ALU_Output[19]
port 39 nsew signal output
rlabel metal3 s 200 356328 800 356448 6 ALU_Output[1]
port 40 nsew signal output
rlabel metal2 s 68282 200 68338 800 6 ALU_Output[20]
port 41 nsew signal output
rlabel metal2 s 110142 379200 110198 379800 6 ALU_Output[21]
port 42 nsew signal output
rlabel metal3 s 194200 74128 194800 74248 6 ALU_Output[22]
port 43 nsew signal output
rlabel metal3 s 200 135328 800 135448 6 ALU_Output[23]
port 44 nsew signal output
rlabel metal3 s 200 144168 800 144288 6 ALU_Output[24]
port 45 nsew signal output
rlabel metal3 s 194200 2048 194800 2168 6 ALU_Output[25]
port 46 nsew signal output
rlabel metal2 s 13542 379200 13598 379800 6 ALU_Output[26]
port 47 nsew signal output
rlabel metal2 s 120446 200 120502 800 6 ALU_Output[27]
port 48 nsew signal output
rlabel metal2 s 94042 379200 94098 379800 6 ALU_Output[28]
port 49 nsew signal output
rlabel metal3 s 194200 252288 194800 252408 6 ALU_Output[29]
port 50 nsew signal output
rlabel metal2 s 61842 379200 61898 379800 6 ALU_Output[2]
port 51 nsew signal output
rlabel metal3 s 200 377408 800 377528 6 ALU_Output[30]
port 52 nsew signal output
rlabel metal3 s 194200 312128 194800 312248 6 ALU_Output[31]
port 53 nsew signal output
rlabel metal3 s 200 348168 800 348288 6 ALU_Output[32]
port 54 nsew signal output
rlabel metal2 s 152646 200 152702 800 6 ALU_Output[33]
port 55 nsew signal output
rlabel metal3 s 200 148248 800 148368 6 ALU_Output[34]
port 56 nsew signal output
rlabel metal3 s 200 309408 800 309528 6 ALU_Output[35]
port 57 nsew signal output
rlabel metal2 s 15474 200 15530 800 6 ALU_Output[36]
port 58 nsew signal output
rlabel metal3 s 200 169328 800 169448 6 ALU_Output[37]
port 59 nsew signal output
rlabel metal3 s 194200 290368 194800 290488 6 ALU_Output[38]
port 60 nsew signal output
rlabel metal2 s 47674 200 47730 800 6 ALU_Output[39]
port 61 nsew signal output
rlabel metal3 s 200 233248 800 233368 6 ALU_Output[3]
port 62 nsew signal output
rlabel metal3 s 194200 99288 194800 99408 6 ALU_Output[40]
port 63 nsew signal output
rlabel metal3 s 194200 358368 194800 358488 6 ALU_Output[41]
port 64 nsew signal output
rlabel metal3 s 194200 91128 194800 91248 6 ALU_Output[42]
port 65 nsew signal output
rlabel metal2 s 63774 200 63830 800 6 ALU_Output[43]
port 66 nsew signal output
rlabel metal3 s 200 301248 800 301368 6 ALU_Output[44]
port 67 nsew signal output
rlabel metal3 s 194200 53048 194800 53168 6 ALU_Output[45]
port 68 nsew signal output
rlabel metal3 s 200 373328 800 373448 6 ALU_Output[46]
port 69 nsew signal output
rlabel metal3 s 194200 137368 194800 137488 6 ALU_Output[47]
port 70 nsew signal output
rlabel metal2 s 74078 379200 74134 379800 6 ALU_Output[48]
port 71 nsew signal output
rlabel metal3 s 194200 159128 194800 159248 6 ALU_Output[49]
port 72 nsew signal output
rlabel metal2 s 21914 379200 21970 379800 6 ALU_Output[4]
port 73 nsew signal output
rlabel metal3 s 200 331168 800 331288 6 ALU_Output[50]
port 74 nsew signal output
rlabel metal3 s 200 335248 800 335368 6 ALU_Output[51]
port 75 nsew signal output
rlabel metal2 s 166814 379200 166870 379800 6 ALU_Output[52]
port 76 nsew signal output
rlabel metal3 s 200 55088 800 55208 6 ALU_Output[53]
port 77 nsew signal output
rlabel metal3 s 194200 133288 194800 133408 6 ALU_Output[54]
port 78 nsew signal output
rlabel metal3 s 194200 367208 194800 367328 6 ALU_Output[55]
port 79 nsew signal output
rlabel metal2 s 194506 379200 194562 379800 6 ALU_Output[56]
port 80 nsew signal output
rlabel metal2 s 31574 200 31630 800 6 ALU_Output[57]
port 81 nsew signal output
rlabel metal2 s 140410 200 140466 800 6 ALU_Output[58]
port 82 nsew signal output
rlabel metal3 s 194200 375368 194800 375488 6 ALU_Output[59]
port 83 nsew signal output
rlabel metal3 s 200 42168 800 42288 6 ALU_Output[5]
port 84 nsew signal output
rlabel metal3 s 200 314168 800 314288 6 ALU_Output[60]
port 85 nsew signal output
rlabel metal2 s 179050 379200 179106 379800 6 ALU_Output[61]
port 86 nsew signal output
rlabel metal2 s 88246 200 88302 800 6 ALU_Output[62]
port 87 nsew signal output
rlabel metal3 s 200 178168 800 178288 6 ALU_Output[63]
port 88 nsew signal output
rlabel metal2 s 84382 200 84438 800 6 ALU_Output[64]
port 89 nsew signal output
rlabel metal3 s 200 59168 800 59288 6 ALU_Output[65]
port 90 nsew signal output
rlabel metal2 s 34150 379200 34206 379800 6 ALU_Output[66]
port 91 nsew signal output
rlabel metal3 s 194200 235288 194800 235408 6 ALU_Output[67]
port 92 nsew signal output
rlabel metal3 s 194200 125128 194800 125248 6 ALU_Output[68]
port 93 nsew signal output
rlabel metal2 s 45742 379200 45798 379800 6 ALU_Output[69]
port 94 nsew signal output
rlabel metal2 s 98550 379200 98606 379800 6 ALU_Output[6]
port 95 nsew signal output
rlabel metal2 s 43810 200 43866 800 6 ALU_Output[70]
port 96 nsew signal output
rlabel metal3 s 194200 265208 194800 265328 6 ALU_Output[71]
port 97 nsew signal output
rlabel metal3 s 200 292408 800 292528 6 ALU_Output[72]
port 98 nsew signal output
rlabel metal3 s 194200 27208 194800 27328 6 ALU_Output[73]
port 99 nsew signal output
rlabel metal2 s 146850 379200 146906 379800 6 ALU_Output[74]
port 100 nsew signal output
rlabel metal2 s 108210 200 108266 800 6 ALU_Output[75]
port 101 nsew signal output
rlabel metal3 s 194200 70048 194800 70168 6 ALU_Output[76]
port 102 nsew signal output
rlabel metal2 s 126242 379200 126298 379800 6 ALU_Output[77]
port 103 nsew signal output
rlabel metal3 s 194200 112208 194800 112328 6 ALU_Output[78]
port 104 nsew signal output
rlabel metal3 s 200 165248 800 165368 6 ALU_Output[79]
port 105 nsew signal output
rlabel metal3 s 200 254328 800 254448 6 ALU_Output[7]
port 106 nsew signal output
rlabel metal2 s 182914 379200 182970 379800 6 ALU_Output[80]
port 107 nsew signal output
rlabel metal3 s 200 365168 800 365288 6 ALU_Output[81]
port 108 nsew signal output
rlabel metal3 s 200 110168 800 110288 6 ALU_Output[82]
port 109 nsew signal output
rlabel metal3 s 200 360408 800 360528 6 ALU_Output[83]
port 110 nsew signal output
rlabel metal2 s 9678 379200 9734 379800 6 ALU_Output[84]
port 111 nsew signal output
rlabel metal2 s 25778 379200 25834 379800 6 ALU_Output[85]
port 112 nsew signal output
rlabel metal3 s 200 16328 800 16448 6 ALU_Output[86]
port 113 nsew signal output
rlabel metal3 s 194200 95208 194800 95328 6 ALU_Output[87]
port 114 nsew signal output
rlabel metal3 s 194200 205368 194800 205488 6 ALU_Output[88]
port 115 nsew signal output
rlabel metal3 s 200 84328 800 84448 6 ALU_Output[89]
port 116 nsew signal output
rlabel metal3 s 194200 248208 194800 248328 6 ALU_Output[8]
port 117 nsew signal output
rlabel metal3 s 200 25168 800 25288 6 ALU_Output[90]
port 118 nsew signal output
rlabel metal3 s 200 369248 800 369368 6 ALU_Output[91]
port 119 nsew signal output
rlabel metal2 s 172610 200 172666 800 6 ALU_Output[92]
port 120 nsew signal output
rlabel metal3 s 194200 269288 194800 269408 6 ALU_Output[93]
port 121 nsew signal output
rlabel metal2 s 36082 200 36138 800 6 ALU_Output[94]
port 122 nsew signal output
rlabel metal3 s 200 140088 800 140208 6 ALU_Output[95]
port 123 nsew signal output
rlabel metal3 s 200 271328 800 271448 6 ALU_Output[96]
port 124 nsew signal output
rlabel metal2 s 29642 379200 29698 379800 6 ALU_Output[97]
port 125 nsew signal output
rlabel metal3 s 194200 180208 194800 180328 6 ALU_Output[98]
port 126 nsew signal output
rlabel metal3 s 194200 333208 194800 333328 6 ALU_Output[99]
port 127 nsew signal output
rlabel metal3 s 194200 176128 194800 176248 6 ALU_Output[9]
port 128 nsew signal output
rlabel metal2 s 100482 200 100538 800 6 Exception[0]
port 129 nsew signal output
rlabel metal3 s 194200 244128 194800 244248 6 Exception[1]
port 130 nsew signal output
rlabel metal3 s 200 152328 800 152448 6 Exception[2]
port 131 nsew signal output
rlabel metal3 s 200 118328 800 118448 6 Exception[3]
port 132 nsew signal output
rlabel metal2 s 156510 200 156566 800 6 Operation[0]
port 133 nsew signal input
rlabel metal3 s 200 50328 800 50448 6 Operation[1]
port 134 nsew signal input
rlabel metal2 s 150714 379200 150770 379800 6 Operation[2]
port 135 nsew signal input
rlabel metal3 s 194200 239368 194800 239488 6 Operation[3]
port 136 nsew signal input
rlabel metal3 s 194200 40128 194800 40248 6 Overflow[0]
port 137 nsew signal output
rlabel metal3 s 200 106088 800 106208 6 Overflow[1]
port 138 nsew signal output
rlabel metal3 s 200 280168 800 280288 6 Overflow[2]
port 139 nsew signal output
rlabel metal3 s 200 237328 800 237448 6 Overflow[3]
port 140 nsew signal output
rlabel metal3 s 200 343408 800 343528 6 Underflow[0]
port 141 nsew signal output
rlabel metal3 s 194200 273368 194800 273488 6 Underflow[1]
port 142 nsew signal output
rlabel metal2 s 168746 200 168802 800 6 Underflow[2]
port 143 nsew signal output
rlabel metal3 s 200 63248 800 63368 6 Underflow[3]
port 144 nsew signal output
rlabel metal2 s 160374 200 160430 800 6 clk
port 145 nsew signal input
rlabel metal3 s 200 305328 800 305448 6 iCE
port 146 nsew signal input
rlabel metal3 s 194200 171368 194800 171488 6 i_operand_sel
port 147 nsew signal input
rlabel metal2 s 86314 379200 86370 379800 6 i_rst
port 148 nsew signal input
rlabel metal2 s 174542 379200 174598 379800 6 operand[0]
port 149 nsew signal input
rlabel metal2 s 90178 379200 90234 379800 6 operand[100]
port 150 nsew signal input
rlabel metal3 s 194200 167288 194800 167408 6 operand[101]
port 151 nsew signal input
rlabel metal3 s 194200 324368 194800 324488 6 operand[102]
port 152 nsew signal input
rlabel metal3 s 194200 142128 194800 142248 6 operand[103]
port 153 nsew signal input
rlabel metal3 s 200 46248 800 46368 6 operand[104]
port 154 nsew signal input
rlabel metal3 s 194200 282208 194800 282328 6 operand[105]
port 155 nsew signal input
rlabel metal3 s 194200 48288 194800 48408 6 operand[106]
port 156 nsew signal input
rlabel metal3 s 194200 354288 194800 354408 6 operand[107]
port 157 nsew signal input
rlabel metal3 s 194200 10208 194800 10328 6 operand[108]
port 158 nsew signal input
rlabel metal2 s 70214 379200 70270 379800 6 operand[109]
port 159 nsew signal input
rlabel metal2 s 27710 200 27766 800 6 operand[10]
port 160 nsew signal input
rlabel metal3 s 194200 146208 194800 146328 6 operand[110]
port 161 nsew signal input
rlabel metal2 s 124310 200 124366 800 6 operand[111]
port 162 nsew signal input
rlabel metal3 s 194200 184288 194800 184408 6 operand[112]
port 163 nsew signal input
rlabel metal3 s 200 93168 800 93288 6 operand[113]
port 164 nsew signal input
rlabel metal3 s 200 203328 800 203448 6 operand[114]
port 165 nsew signal input
rlabel metal2 s 134614 379200 134670 379800 6 operand[115]
port 166 nsew signal input
rlabel metal3 s 194200 307368 194800 307488 6 operand[116]
port 167 nsew signal input
rlabel metal3 s 194200 218288 194800 218408 6 operand[117]
port 168 nsew signal input
rlabel metal3 s 200 72088 800 72208 6 operand[118]
port 169 nsew signal input
rlabel metal2 s 138478 379200 138534 379800 6 operand[119]
port 170 nsew signal input
rlabel metal3 s 200 191088 800 191208 6 operand[11]
port 171 nsew signal input
rlabel metal3 s 200 29248 800 29368 6 operand[120]
port 172 nsew signal input
rlabel metal3 s 200 101328 800 101448 6 operand[121]
port 173 nsew signal input
rlabel metal3 s 200 288328 800 288448 6 operand[122]
port 174 nsew signal input
rlabel metal2 s 158442 379200 158498 379800 6 operand[123]
port 175 nsew signal input
rlabel metal2 s 66350 379200 66406 379800 6 operand[124]
port 176 nsew signal input
rlabel metal3 s 200 161168 800 161288 6 operand[125]
port 177 nsew signal input
rlabel metal3 s 200 182248 800 182368 6 operand[126]
port 178 nsew signal input
rlabel metal3 s 194200 222368 194800 222488 6 operand[127]
port 179 nsew signal input
rlabel metal3 s 194200 210128 194800 210248 6 operand[12]
port 180 nsew signal input
rlabel metal3 s 200 76168 800 76288 6 operand[13]
port 181 nsew signal input
rlabel metal3 s 194200 193128 194800 193248 6 operand[14]
port 182 nsew signal input
rlabel metal3 s 194200 120368 194800 120488 6 operand[15]
port 183 nsew signal input
rlabel metal3 s 194200 36048 194800 36168 6 operand[16]
port 184 nsew signal input
rlabel metal3 s 200 195168 800 195288 6 operand[17]
port 185 nsew signal input
rlabel metal3 s 194200 316208 194800 316328 6 operand[18]
port 186 nsew signal input
rlabel metal2 s 136546 200 136602 800 6 operand[19]
port 187 nsew signal input
rlabel metal2 s 192574 200 192630 800 6 operand[1]
port 188 nsew signal input
rlabel metal3 s 194200 103368 194800 103488 6 operand[20]
port 189 nsew signal input
rlabel metal2 s 57978 379200 58034 379800 6 operand[21]
port 190 nsew signal input
rlabel metal2 s 132682 200 132738 800 6 operand[22]
port 191 nsew signal input
rlabel metal2 s 23846 200 23902 800 6 operand[23]
port 192 nsew signal input
rlabel metal3 s 200 33328 800 33448 6 operand[24]
port 193 nsew signal input
rlabel metal3 s 194200 201288 194800 201408 6 operand[25]
port 194 nsew signal input
rlabel metal3 s 194200 295128 194800 295248 6 operand[26]
port 195 nsew signal input
rlabel metal2 s 92110 200 92166 800 6 operand[27]
port 196 nsew signal input
rlabel metal3 s 194200 363128 194800 363248 6 operand[28]
port 197 nsew signal input
rlabel metal3 s 200 12248 800 12368 6 operand[29]
port 198 nsew signal input
rlabel metal2 s 188710 200 188766 800 6 operand[2]
port 199 nsew signal input
rlabel metal3 s 194200 371288 194800 371408 6 operand[30]
port 200 nsew signal input
rlabel metal2 s 184846 200 184902 800 6 operand[31]
port 201 nsew signal input
rlabel metal2 s 76010 200 76066 800 6 operand[32]
port 202 nsew signal input
rlabel metal2 s 11610 200 11666 800 6 operand[33]
port 203 nsew signal input
rlabel metal3 s 194200 57128 194800 57248 6 operand[34]
port 204 nsew signal input
rlabel metal3 s 194200 129208 194800 129328 6 operand[35]
port 205 nsew signal input
rlabel metal2 s 82450 379200 82506 379800 6 operand[36]
port 206 nsew signal input
rlabel metal3 s 194200 286288 194800 286408 6 operand[37]
port 207 nsew signal input
rlabel metal3 s 200 322328 800 322448 6 operand[38]
port 208 nsew signal input
rlabel metal3 s 200 339328 800 339448 6 operand[39]
port 209 nsew signal input
rlabel metal3 s 200 21088 800 21208 6 operand[3]
port 210 nsew signal input
rlabel metal2 s 7746 200 7802 800 6 operand[40]
port 211 nsew signal input
rlabel metal2 s 52182 200 52238 800 6 operand[41]
port 212 nsew signal input
rlabel metal3 s 194200 197208 194800 197328 6 operand[42]
port 213 nsew signal input
rlabel metal2 s 144274 200 144330 800 6 operand[43]
port 214 nsew signal input
rlabel metal2 s 162950 379200 163006 379800 6 operand[44]
port 215 nsew signal input
rlabel metal3 s 194200 350208 194800 350328 6 operand[45]
port 216 nsew signal input
rlabel metal2 s 1950 379200 2006 379800 6 operand[46]
port 217 nsew signal input
rlabel metal3 s 200 186328 800 186448 6 operand[47]
port 218 nsew signal input
rlabel metal3 s 194200 227128 194800 227248 6 operand[48]
port 219 nsew signal input
rlabel metal3 s 194200 346128 194800 346248 6 operand[49]
port 220 nsew signal input
rlabel metal3 s 200 250248 800 250368 6 operand[4]
port 221 nsew signal input
rlabel metal3 s 194200 278128 194800 278248 6 operand[50]
port 222 nsew signal input
rlabel metal3 s 194200 154368 194800 154488 6 operand[51]
port 223 nsew signal input
rlabel metal2 s 176474 200 176530 800 6 operand[52]
port 224 nsew signal input
rlabel metal2 s 190642 379200 190698 379800 6 operand[53]
port 225 nsew signal input
rlabel metal2 s 38014 379200 38070 379800 6 operand[54]
port 226 nsew signal input
rlabel metal2 s 79874 200 79930 800 6 operand[55]
port 227 nsew signal input
rlabel metal3 s 200 157088 800 157208 6 operand[56]
port 228 nsew signal input
rlabel metal3 s 200 114248 800 114368 6 operand[57]
port 229 nsew signal input
rlabel metal3 s 194200 150288 194800 150408 6 operand[58]
port 230 nsew signal input
rlabel metal3 s 200 220328 800 220448 6 operand[59]
port 231 nsew signal input
rlabel metal3 s 194200 78208 194800 78328 6 operand[5]
port 232 nsew signal input
rlabel metal2 s 39946 200 40002 800 6 operand[60]
port 233 nsew signal input
rlabel metal2 s 128174 200 128230 800 6 operand[61]
port 234 nsew signal input
rlabel metal3 s 194200 188368 194800 188488 6 operand[62]
port 235 nsew signal input
rlabel metal2 s 170678 379200 170734 379800 6 operand[63]
port 236 nsew signal input
rlabel metal3 s 194200 320288 194800 320408 6 operand[64]
port 237 nsew signal input
rlabel metal3 s 194200 87048 194800 87168 6 operand[65]
port 238 nsew signal input
rlabel metal3 s 200 89088 800 89208 6 operand[66]
port 239 nsew signal input
rlabel metal3 s 200 4088 800 4208 6 operand[67]
port 240 nsew signal input
rlabel metal2 s 3882 200 3938 800 6 operand[68]
port 241 nsew signal input
rlabel metal3 s 194200 329128 194800 329248 6 operand[69]
port 242 nsew signal input
rlabel metal2 s 154578 379200 154634 379800 6 operand[6]
port 243 nsew signal input
rlabel metal3 s 194200 108128 194800 108248 6 operand[70]
port 244 nsew signal input
rlabel metal2 s 142342 379200 142398 379800 6 operand[71]
port 245 nsew signal input
rlabel metal3 s 200 123088 800 123208 6 operand[72]
port 246 nsew signal input
rlabel metal3 s 200 131248 800 131368 6 operand[73]
port 247 nsew signal input
rlabel metal2 s 180982 200 181038 800 6 operand[74]
port 248 nsew signal input
rlabel metal2 s 18 200 74 800 6 operand[75]
port 249 nsew signal input
rlabel metal3 s 194200 19048 194800 19168 6 operand[76]
port 250 nsew signal input
rlabel metal3 s 200 174088 800 174208 6 operand[77]
port 251 nsew signal input
rlabel metal3 s 200 284248 800 284368 6 operand[78]
port 252 nsew signal input
rlabel metal3 s 200 80248 800 80368 6 operand[79]
port 253 nsew signal input
rlabel metal3 s 200 127168 800 127288 6 operand[7]
port 254 nsew signal input
rlabel metal2 s 56046 200 56102 800 6 operand[80]
port 255 nsew signal input
rlabel metal2 s 19982 200 20038 800 6 operand[81]
port 256 nsew signal input
rlabel metal2 s 77942 379200 77998 379800 6 operand[82]
port 257 nsew signal input
rlabel metal2 s 18050 379200 18106 379800 6 operand[83]
port 258 nsew signal input
rlabel metal2 s 148782 200 148838 800 6 operand[84]
port 259 nsew signal input
rlabel metal2 s 122378 379200 122434 379800 6 operand[85]
port 260 nsew signal input
rlabel metal3 s 194200 163208 194800 163328 6 operand[86]
port 261 nsew signal input
rlabel metal3 s 200 212168 800 212288 6 operand[87]
port 262 nsew signal input
rlabel metal3 s 194200 303288 194800 303408 6 operand[88]
port 263 nsew signal input
rlabel metal2 s 59910 200 59966 800 6 operand[89]
port 264 nsew signal input
rlabel metal2 s 104346 200 104402 800 6 operand[8]
port 265 nsew signal input
rlabel metal3 s 200 38088 800 38208 6 operand[90]
port 266 nsew signal input
rlabel metal3 s 194200 299208 194800 299328 6 operand[91]
port 267 nsew signal input
rlabel metal2 s 164882 200 164938 800 6 operand[92]
port 268 nsew signal input
rlabel metal2 s 106278 379200 106334 379800 6 operand[93]
port 269 nsew signal input
rlabel metal2 s 102414 379200 102470 379800 6 operand[94]
port 270 nsew signal input
rlabel metal3 s 200 276088 800 276208 6 operand[95]
port 271 nsew signal input
rlabel metal3 s 200 326408 800 326528 6 operand[96]
port 272 nsew signal input
rlabel metal3 s 194200 6128 194800 6248 6 operand[97]
port 273 nsew signal input
rlabel metal3 s 200 67328 800 67448 6 operand[98]
port 274 nsew signal input
rlabel metal3 s 200 242088 800 242208 6 operand[99]
port 275 nsew signal input
rlabel metal3 s 194200 231208 194800 231328 6 operand[9]
port 276 nsew signal input
rlabel metal4 s 4208 2128 4528 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 377584 6 vccd1
port 277 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 377584 6 vssd1
port 278 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 377584 6 vssd1
port 278 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 377584 6 vssd1
port 278 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 377584 6 vssd1
port 278 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 377584 6 vssd1
port 278 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 377584 6 vssd1
port 278 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 195000 380000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 176177958
string GDS_FILE /home/baungarten/Caravel_4_ALU_fixed/openlane/ALL_ALU/runs/23_02_20_07_27/results/signoff/Top_Module_4_ALU.magic.gds
string GDS_START 1647468
<< end >>

