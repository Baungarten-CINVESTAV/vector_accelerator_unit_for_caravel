* NGSPICE file created from ALU.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

.subckt ALU ALU_Output[0] ALU_Output[10] ALU_Output[11] ALU_Output[12] ALU_Output[13]
+ ALU_Output[14] ALU_Output[15] ALU_Output[16] ALU_Output[17] ALU_Output[18] ALU_Output[19]
+ ALU_Output[1] ALU_Output[20] ALU_Output[21] ALU_Output[22] ALU_Output[23] ALU_Output[24]
+ ALU_Output[25] ALU_Output[26] ALU_Output[27] ALU_Output[28] ALU_Output[29] ALU_Output[2]
+ ALU_Output[30] ALU_Output[31] ALU_Output[3] ALU_Output[4] ALU_Output[5] ALU_Output[6]
+ ALU_Output[7] ALU_Output[8] ALU_Output[9] Exception Operation[0] Operation[1] Operation[2]
+ Operation[3] Overflow Underflow a_operand[0] a_operand[10] a_operand[11] a_operand[12]
+ a_operand[13] a_operand[14] a_operand[15] a_operand[16] a_operand[17] a_operand[18]
+ a_operand[19] a_operand[1] a_operand[20] a_operand[21] a_operand[22] a_operand[23]
+ a_operand[24] a_operand[25] a_operand[26] a_operand[27] a_operand[28] a_operand[29]
+ a_operand[2] a_operand[30] a_operand[31] a_operand[3] a_operand[4] a_operand[5]
+ a_operand[6] a_operand[7] a_operand[8] a_operand[9] b_operand[0] b_operand[10] b_operand[11]
+ b_operand[12] b_operand[13] b_operand[14] b_operand[15] b_operand[16] b_operand[17]
+ b_operand[18] b_operand[19] b_operand[1] b_operand[20] b_operand[21] b_operand[22]
+ b_operand[23] b_operand[24] b_operand[25] b_operand[26] b_operand[27] b_operand[28]
+ b_operand[29] b_operand[2] b_operand[30] b_operand[31] b_operand[3] b_operand[4]
+ b_operand[5] b_operand[6] b_operand[7] b_operand[8] b_operand[9] vccd1 vssd1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12222__C _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4777_ MuI._0312_ MuI._0313_ MuI._0323_ vssd1 vssd1 vccd1 vccd1 MuI._0498_ sky130_fd_sc_hd__nor3_1
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ _02309_ _02310_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__nor3_1
X_06883_ _04165_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__buf_4
XFILLER_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6516_ MuI._2409_ MuI._2410_ vssd1 vssd1 vccd1 vccd1 MuI._2411_ sky130_fd_sc_hd__or2_1
XMuI._3728_ MuI._2825_ MuI._2827_ vssd1 vssd1 vccd1 vccd1 MuI._2828_ sky130_fd_sc_hd__nor2_1
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08622_ _01237_ _01239_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__and2_1
XFILLER_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6447_ MuI._2331_ MuI._2334_ vssd1 vssd1 vccd1 vccd1 MuI._2335_ sky130_fd_sc_hd__and2b_1
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3659_ MuI.a_operand\[15\] vssd1 vssd1 vccd1 vccd1 MuI._2605_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07613__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _01164_ _01168_ _01170_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__o21ba_1
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6378_ MuI._2826_ MuI._0603_ MuI._2594_ MuI._2797_ vssd1 vssd1 vccd1 vccd1 MuI._2259_
+ sky130_fd_sc_hd__and4_1
X_07504_ _00107_ _00108_ _00120_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4209__B1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__B2 _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07332__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ _01099_ _01101_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__nor2_2
XFILLER_196_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5329_ MuI._0969_ MuI._0970_ MuI._0971_ vssd1 vssd1 vccd1 vccd1 MuI._1105_ sky130_fd_sc_hd__and3_1
XFILLER_168_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _00037_ _00043_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__nor2_1
XFILLER_196_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4091__C MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07366_ _06565_ _02485_ _06476_ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nand4_1
XFILLER_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11397__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _01720_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__and2_1
XFILLER_176_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07297_ net40 vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__clkbuf_4
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09036_ _01204_ _01208_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__nor2_1
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06899__A _04338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__A2 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _02599_ _02088_ _02598_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__or3b_1
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12132__C _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _02490_ _02491_ _02517_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07226__C net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _03525_ _06613_ _04558_ _04557_ _04918_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__a32o_1
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _02720_ _02805_ _02730_ AuI.result\[20\] vssd1 vssd1 vccd1 vccd1 _05765_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5659__A MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _02871_ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5660__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__B1 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3671__A1 MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07828__A2 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _06429_ _04725_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__nand2_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10713_ _03429_ _03430_ _03431_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__a21o_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ _02571_ _04159_ _04348_ _04357_ _04490_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__o311a_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ FuI.Integer\[29\] _06045_ _02717_ _05917_ vssd1 vssd1 vccd1 vccd1 _06347_
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _03389_ _02984_ _00036_ _00059_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand4_1
XFILLER_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__A1 _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09169__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ _03108_ _03111_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nand2_1
X_13363_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__inv_2
XANTENNA__10596__B1 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09805__A2_N net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _05149_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13294_ _06146_ _06151_ _02833_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21ai_1
XFILLER_182_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _03525_ _04983_ _04944_ _04943_ _05123_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a32o_2
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1623_ AuI._0259_ AuI._0789_ AuI._0790_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[18\]
+ sky130_fd_sc_hd__o211a_1
X_12176_ _04800_ _02941_ _02938_ AuI.result\[13\] vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4700_ MuI._0266_ MuI._0272_ vssd1 vssd1 vccd1 vccd1 MuI._0413_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12323__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5680_ MuI._1487_ MuI._1488_ MuI._1489_ vssd1 vssd1 vccd1 vccd1 MuI._1491_ sky130_fd_sc_hd__a21o_1
XFILLER_150_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1554_ AuI._0701_ AuI._0728_ AuI._0733_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0734_
+ sky130_fd_sc_hd__o22a_1
X_11127_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__xnor2_4
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._560_ AuI.pe._074_ AuI.pe._109_ AuI.pe._111_ AuI.pe._116_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[9\] sky130_fd_sc_hd__o22a_1
XMuI._4631_ MuI._0212_ MuI._0211_ vssd1 vssd1 vccd1 vccd1 MuI._0337_ sky130_fd_sc_hd__nor2_1
XFILLER_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11848__B1 _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _03803_ _03804_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__xor2_2
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1485_ AuI._0524_ AuI._0527_ vssd1 vssd1 vccd1 vccd1 AuI._0671_ sky130_fd_sc_hd__nor2_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07516__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._491_ AuI.pe._386_ AuI.pe._000_ AuI.pe._384_ vssd1 vssd1 vccd1 vccd1 AuI.pe._053_
+ sky130_fd_sc_hd__and3_2
XANTENNA__11312__A2 _04076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4562_ MuI._0254_ MuI._0260_ vssd1 vssd1 vccd1 vccd1 MuI._0261_ sky130_fd_sc_hd__xor2_1
X_10009_ _02665_ _02666_ _02676_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__nand3_1
XFILLER_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__B _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6301_ MuI._0889_ MuI._1494_ MuI._2172_ vssd1 vssd1 vccd1 vccd1 MuI._2174_ sky130_fd_sc_hd__a21oi_1
XMuI._3513_ MuI._0394_ MuI._0548_ MuI._0988_ vssd1 vssd1 vccd1 vccd1 MuI._0999_ sky130_fd_sc_hd__nor3_2
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08529__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4493_ MuI._2975_ MuI._2451_ MuI._2845_ MuI._2440_ vssd1 vssd1 vccd1 vccd1 MuI._0186_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6232_ MuI._2092_ MuI._2097_ vssd1 vssd1 vccd1 vccd1 MuI._2098_ sky130_fd_sc_hd__xnor2_1
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3444_ MuI._0196_ MuI._0218_ MuI._0229_ vssd1 vssd1 vccd1 vccd1 MuI._0240_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07152__B _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12993__B _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6163_ MuI._2019_ MuI._2020_ MuI._2021_ vssd1 vssd1 vccd1 vccd1 MuI._2023_ sky130_fd_sc_hd__or3_1
XFILLER_177_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4623__D MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__A _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5114_ MuI._0866_ MuI._0868_ vssd1 vssd1 vccd1 vccd1 MuI._0869_ sky130_fd_sc_hd__nor2_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _06516_ _06517_ _06518_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__a22oi_1
XMuI._6094_ MuI._1942_ MuI._1946_ vssd1 vssd1 vccd1 vccd1 MuI._1947_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5045_ MuI._0283_ MuI._0786_ MuI._0789_ MuI._0792_ vssd1 vssd1 vccd1 vccd1 MuI._0793_
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__11379__A2 _04000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__C1 _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07151_ _06450_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__nor2_2
XFILLER_158_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _06295_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08711__B _01325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5947_ MuI._1738_ MuI._1739_ vssd1 vssd1 vccd1 vccd1 MuI._1785_ sky130_fd_sc_hd__nand2_1
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13329__B _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout105 FuI.a_operand\[30\] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._827_ AuI.operand_a\[27\] AuI.pe._273_ AuI.operand_a\[28\] vssd1 vssd1 vccd1
+ vccd1 AuI.pe._364_ sky130_fd_sc_hd__a21o_1
Xfanout116 net48 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_4
XFILLER_141_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout127 net27 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_2
XFILLER_86_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5878_ MuI._1707_ MuI._1708_ vssd1 vssd1 vccd1 vccd1 MuI._1709_ sky130_fd_sc_hd__nand2_1
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07984_ _00600_ _00601_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__and2b_1
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4142__A2 MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4829_ MuI._0552_ MuI._0553_ MuI._0554_ vssd1 vssd1 vccd1 vccd1 MuI._0555_ sky130_fd_sc_hd__or3_1
XAuI.pe._758_ AuI.pe.significand\[5\] AuI.pe._213_ AuI.pe._078_ AuI.pe._201_ AuI.pe._301_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._302_ sky130_fd_sc_hd__a221o_1
X_09723_ _02280_ _02279_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__nor2_1
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11839__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06935_ _04725_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__buf_4
XANTENNA__11303__A2 _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4086__C MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12500__A1 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._689_ AuI.pe._106_ AuI.pe._112_ AuI.pe._230_ AuI.pe._231_ AuI.pe._236_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._237_ sky130_fd_sc_hd__a2111o_1
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _02247_ _02245_ _02246_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__nand3_1
XFILLER_95_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06866_ _03982_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07343__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _01220_ _01221_ _01222_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__o21bai_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06797_ _03239_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__and3_1
X_09585_ _02334_ _00266_ _04294_ _01332_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a22o_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1308__A0 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._496__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _01152_ _01142_ _01151_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__nand3_1
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13461__C1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4533__D MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _06601_ _00085_ _04585_ _06606_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__a22oi_1
XFILLER_211_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07418_ _00035_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__buf_4
XANTENNA_AuI.pe._620__D AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ _01007_ _01008_ _01014_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__and3_1
XFILLER_211_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3727__A MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _06646_ _06648_ _06647_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__a21o_1
XFILLER_192_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _06593_ _06477_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__and2_1
XFILLER_191_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09019_ _01237_ _01239_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__xnor2_1
X_10291_ _03432_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__buf_4
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12030_ _04849_ _04850_ _04830_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09735__A2 _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6195__D MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12932_ _05803_ _05819_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xnor2_1
XAuI._1270_ AuI._0460_ AuI._0470_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[11\]
+ sky130_fd_sc_hd__xnor2_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08349__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _05661_ _05663_ _05745_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__or3_1
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11814_ _06428_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__nor2_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _02628_ _05576_ _02596_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a21o_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09120__B1 _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _04544_ _04525_ _04526_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__nand3_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6712__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5836__B MuI._1662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _04469_ _04470_ _04428_ _04429_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a211o_1
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3637__A MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13415_ _06289_ _06292_ _06327_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or3_1
XFuI._148__154 vssd1 vssd1 vccd1 vccd1 FuI._148__154/HI net154 sky130_fd_sc_hd__conb_1
X_10627_ _03615_ _04369_ _04456_ _03550_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__a22oi_1
XFILLER_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09423__A1 _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09423__B2 _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5149__B2 MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10033__A2 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13346_ _05700_ _06205_ _02830_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08234__D _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10558_ _03091_ _03093_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__nand2_1
XAuI._0985_ AuI._0193_ AuI._0196_ vssd1 vssd1 vccd1 vccd1 AuI._0197_ sky130_fd_sc_hd__nor2_1
XANTENNA__08812__A _01391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0825__A2 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6850_ MuI._2678_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[18\] sky130_fd_sc_hd__nor2_1
XFILLER_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13277_ _06106_ _06124_ _06105_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__a21bo_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10489_ _03191_ _03189_ _03190_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__nand3_1
XANTENNA__08531__B _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5801_ MuI._1607_ MuI._1622_ MuI._1623_ vssd1 vssd1 vccd1 vccd1 MuI._1624_ sky130_fd_sc_hd__and3_1
XFILLER_142_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4372__A2 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6781_ MuI._2685_ MuI._2591_ vssd1 vssd1 vccd1 vccd1 MuI._2702_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07428__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3993_ MuI._2473_ MuI._2682_ vssd1 vssd1 vccd1 vccd1 MuI._3093_ sky130_fd_sc_hd__nand2_1
XFILLER_97_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12228_ _05063_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4468__A MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5732_ MuI._1545_ MuI._1546_ MuI._1478_ vssd1 vssd1 vccd1 vccd1 MuI._1548_ sky130_fd_sc_hd__a21o_1
XANTENNA__10339__B1_N _00735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6386__C MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__A1 _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1606_ AuI._0710_ AuI._0776_ vssd1 vssd1 vccd1 vccd1 AuI._0777_ sky130_fd_sc_hd__nand2_1
XANTENNA__12730__B2 _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _04904_ _04862_ _04989_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a211oi_4
XAuI.pe._612_ AuI.pe._063_ AuI.pe._097_ AuI.pe._119_ AuI.pe._045_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._165_ sky130_fd_sc_hd__a22o_1
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5663_ MuI._0986_ MuI._1471_ vssd1 vssd1 vccd1 vccd1 MuI._1473_ sky130_fd_sc_hd__nand2_1
XAuI._1537_ AuI._0701_ AuI._0716_ AuI._0718_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0720_
+ sky130_fd_sc_hd__o22a_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4614_ MuI._0112_ MuI._0316_ MuI._0318_ vssd1 vssd1 vccd1 vccd1 MuI._0319_ sky130_fd_sc_hd__a21bo_1
XAuI.pe._543_ AuI.pe.significand\[8\] AuI.pe._375_ AuI.pe._049_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._101_ sky130_fd_sc_hd__or3_4
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5594_ MuI._1393_ MuI._1394_ MuI._1396_ vssd1 vssd1 vccd1 vccd1 MuI._1397_ sky130_fd_sc_hd__nor3b_1
X_06720_ net107 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__clkbuf_8
XFILLER_77_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1468_ AuI._0140_ AuI._0252_ AuI._0610_ AuI._0609_ vssd1 vssd1 vccd1 vccd1 AuI._0654_
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08259__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._474_ AuI.pe._013_ AuI.pe._014_ AuI.pe.significand\[2\] vssd1 vssd1 vccd1
+ vccd1 AuI.pe._038_ sky130_fd_sc_hd__or3_1
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4545_ MuI._0241_ MuI._0242_ vssd1 vssd1 vccd1 vccd1 MuI._0243_ sky130_fd_sc_hd__nor2_1
XFILLER_25_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13038__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1399_ AuI._0587_ AuI._0588_ vssd1 vssd1 vccd1 vccd1 AuI._0589_ sky130_fd_sc_hd__or2b_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4476_ MuI._0164_ MuI._0166_ vssd1 vssd1 vccd1 vccd1 MuI._0167_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09370_ _02420_ _00592_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nand2_2
XMuI._6215_ MuI._2038_ MuI._2078_ MuI._2079_ vssd1 vssd1 vccd1 vccd1 MuI._2080_ sky130_fd_sc_hd__a21o_1
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3427_ MuI.a_operand\[23\] MuI._0032_ MuI._0043_ vssd1 vssd1 vccd1 vccd1 MuI._0054_
+ sky130_fd_sc_hd__and3_1
X_08321_ _00900_ _00937_ _00938_ _00618_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__o211a_1
XFILLER_178_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6146_ MuI._2002_ MuI._2003_ vssd1 vssd1 vccd1 vccd1 MuI._2004_ sky130_fd_sc_hd__nor2_1
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08252_ _00848_ _00847_ _00846_ _00835_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__o211ai_1
XFILLER_178_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__B1 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07203_ net109 vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__buf_4
XMuI._6077_ MuI._1851_ MuI._1859_ vssd1 vssd1 vccd1 vccd1 MuI._1928_ sky130_fd_sc_hd__nand2_1
XFILLER_165_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11132__B _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08183_ _00770_ _00800_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5465__C MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout125_A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13210__A2 _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5028_ MuI._0740_ MuI._0773_ vssd1 vssd1 vccd1 vccd1 MuI._0774_ sky130_fd_sc_hd__nor2_1
X_07134_ _03604_ _04035_ _06433_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a22oi_1
XFILLER_119_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11559__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A2 _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07065_ _06119_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_173_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07728__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07728__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _00563_ _00562_ _00561_ _00545_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__o211a_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09706_ _06504_ _04165_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__and2_1
XFILLER_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06918_ _04542_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__and3_1
XANTENNA__09272__B _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ _00514_ _00504_ _06450_ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__or3_1
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _02228_ _02275_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10849__D _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06849_ _03798_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4544__C MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _02195_ _02196_ _02200_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a21o_1
XFILLER_43_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08519_ _01114_ _01116_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__nor2_1
XFILLER_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _01978_ _01977_ _01970_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a21o_1
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _03660_ _03833_ _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__and3b_1
XANTENNA__07664__B1 _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._154_ net104 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[24\] sky130_fd_sc_hd__clkbuf_1
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3457__A MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__B _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _03909_ _03910_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__nor2_1
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._085_ FuI.a_operand\[23\] FuI._048_ vssd1 vssd1 vccd1 vccd1 FuI._049_ sky130_fd_sc_hd__and2_1
X_13200_ _06105_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and2_1
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10412_ _00712_ _00806_ _03109_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07416__B1 _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11392_ _04391_ _02728_ _04162_ _03494_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_109_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__B _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08632__A _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3607__D MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _03809_ _05595_ _06031_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21o_1
XFILLER_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10343_ _03026_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07248__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _06442_ _00301_ _00259_ _03550_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a22oi_1
X_13062_ _05957_ _05958_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input55_A b_operand[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12712__A1 _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _00270_ _06561_ _04679_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a31o_1
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6500__B1 MuI._1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0852__A2_N net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13268__A2 _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._1322_ net11 net120 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0519_ sky130_fd_sc_hd__mux2_2
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08079__A _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12915_ _05800_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1253_ AuI._0437_ AuI._0452_ AuI._0453_ AuI._0454_ vssd1 vssd1 vccd1 vccd1 AuI._0455_
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4330_ MuI._3292_ MuI._3293_ vssd1 vssd1 vccd1 vccd1 MuI._0007_ sky130_fd_sc_hd__nor2_1
XFILLER_207_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _03798_ _05327_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nand2_1
XFILLER_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1184_ AuI._0307_ AuI._0203_ vssd1 vssd1 vccd1 vccd1 AuI._0390_ sky130_fd_sc_hd__and2_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5269__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4261_ MuI.b_operand\[20\] MuI._2830_ vssd1 vssd1 vccd1 vccd1 MuI._3361_ sky130_fd_sc_hd__nand2_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6000_ MuI._3121_ MuI._3123_ vssd1 vssd1 vccd1 vccd1 MuI._1843_ sky130_fd_sc_hd__nor2_1
X_12777_ _05553_ _05653_ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and3_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13440__A2 _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__B _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4192_ MuI._3290_ MuI._3291_ vssd1 vssd1 vccd1 vccd1 MuI._3292_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _01146_ _06561_ _03047_ _01147_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a22oi_2
XFILLER_30_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10494__D _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _02987_ _04918_ _04450_ _04451_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__nand4_1
XANTENNA__11203__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11203__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _03820_ _05788_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__nand2_1
XANTENNA__09357__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0968_ AuI._0164_ AuI._0169_ AuI._0179_ vssd1 vssd1 vccd1 vccd1 AuI._0180_ sky130_fd_sc_hd__and3_1
XANTENNA__08261__B _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6833_ MuI._2722_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2749_ sky130_fd_sc_hd__and2b_1
XANTENNA__07158__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0899_ AuI._0111_ AuI._0114_ AuI._0117_ AuI._0118_ vssd1 vssd1 vccd1 vccd1 AuI._0119_
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3976_ MuI._3039_ MuI._3059_ vssd1 vssd1 vccd1 vccd1 MuI._3076_ sky130_fd_sc_hd__xnor2_1
XMuI._6764_ MuI._2683_ MuI._2621_ MuI._2626_ vssd1 vssd1 vccd1 vccd1 MuI._2684_ sky130_fd_sc_hd__a21oi_1
X_08870_ _06500_ _06580_ _05025_ _06501_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a22oi_1
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06997__A _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07308__D _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5715_ MuI._1526_ MuI._1528_ MuI._1529_ vssd1 vssd1 vccd1 vccd1 MuI._1530_ sky130_fd_sc_hd__or3_1
XMuI._6695_ MuI._2604_ MuI._2607_ MuI._2505_ vssd1 vssd1 vccd1 vccd1 MuI._2608_ sky130_fd_sc_hd__mux2_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07821_ _00437_ _00436_ _00372_ _00186_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__a211o_1
XFILLER_111_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09804__C _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5646_ MuI._1372_ MuI._1452_ MuI._1453_ vssd1 vssd1 vccd1 vccd1 MuI._1454_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07752_ _00255_ _00256_ _00368_ _00369_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__nand4_2
XAuI.pe._526_ AuI.pe._084_ AuI.pe._070_ vssd1 vssd1 vccd1 vccd1 AuI.pe._085_ sky130_fd_sc_hd__xor2_1
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5577_ MuI._1356_ MuI._1355_ MuI._1347_ vssd1 vssd1 vccd1 vccd1 MuI._1378_ sky130_fd_sc_hd__a21o_1
X_06703_ _02227_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[1\] sky130_fd_sc_hd__clkbuf_4
XFILLER_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07683_ _00267_ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__buf_4
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4528_ MuI._0087_ MuI._0090_ MuI._0091_ vssd1 vssd1 vccd1 vccd1 MuI._0224_ sky130_fd_sc_hd__or3_1
XAuI.pe._457_ AuI.pe._006_ vssd1 vssd1 vccd1 vccd1 AuI.pe._022_ sky130_fd_sc_hd__buf_2
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09422_ _06479_ _06480_ net34 _00082_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__and4_1
XFILLER_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__A2 _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__D _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10966__B _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4588__A1_N MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4459_ MuI._0143_ MuI._0140_ vssd1 vssd1 vccd1 vccd1 MuI._0148_ sky130_fd_sc_hd__xor2_1
XANTENNA__07621__A _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5757__A MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _01933_ _01931_ _01932_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__or3_1
XFILLER_178_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13431__A2 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08304_ _03110_ _00301_ _00259_ _00921_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a22oi_4
X_09284_ _01899_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__nor2_1
XMuI._6129_ MuI._1924_ MuI._1984_ vssd1 vssd1 vccd1 vccd1 MuI._1985_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ net122 _04778_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__nand2_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08166_ _00162_ _05756_ _00783_ _00164_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__a22oi_1
XFILLER_193_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07949__A1 _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07949__B2 _00555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07117_ _06422_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[27\] sky130_fd_sc_hd__clkbuf_1
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _00062_ _06591_ _06584_ _00049_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__a22o_1
XFILLER_161_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07068__A _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ net29 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._6100__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10206__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06700__A _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _01508_ _01509_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__B1 _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09433__D _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5049__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__C net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10961_ _04596_ _03698_ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12700_ _02613_ _05386_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nand2_1
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _03624_ _03623_ _03622_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a21bo_1
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12631_ _02801_ _02875_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__or3_1
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _03733_ _05123_ _05298_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__nand3_1
XFILLER_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11513_ _04250_ _04252_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__and4_1
XFILLER_200_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ _05238_ _05239_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__nor2_1
XFILLER_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._137_ FuI._021_ net143 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[8\] sky130_fd_sc_hd__dlxtn_1
XANTENNA__13186__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__A _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11444_ _04218_ _04219_ _04045_ _04048_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__o211a_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08362__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._068_ FuI.a_operand\[26\] vssd1 vssd1 vccd1 vccd1 FuI._036_ sky130_fd_sc_hd__inv_2
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0822_ AuI._0039_ net14 vssd1 vssd1 vccd1 vccd1 AuI._0042_ sky130_fd_sc_hd__or2_1
X_11375_ _03861_ _03995_ _03994_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__a21oi_2
XFILLER_153_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6721__A0 MuI._2629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ _05966_ _05968_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__or2b_1
XFILLER_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10326_ _00721_ _00720_ _00719_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a21bo_1
XFILLER_180_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._444__A_N AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3830_ MuI._1307_ MuI._1802_ MuI._2440_ vssd1 vssd1 vccd1 vccd1 MuI._2930_ sky130_fd_sc_hd__and3_1
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _03400_ _05981_ _05869_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__a21o_1
X_10257_ _02706_ _02729_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__and2b_1
XFILLER_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3761_ MuI._2860_ MuI._2594_ vssd1 vssd1 vccd1 vccd1 MuI._2861_ sky130_fd_sc_hd__nand2_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _04671_ _02723_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__and2b_1
XFILLER_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5500_ MuI._1282_ MuI._1283_ MuI._1276_ vssd1 vssd1 vccd1 vccd1 MuI._1293_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5827__A2 MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6480_ MuI._2368_ MuI._2370_ vssd1 vssd1 vccd1 vccd1 MuI._2371_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._3650__A MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1042__A AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3692_ MuI._2517_ MuI._2789_ MuI._2791_ MuI._1318_ vssd1 vssd1 vccd1 vccd1 MuI._2792_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5431_ MuI._1202_ MuI._1214_ MuI._1215_ MuI._1216_ vssd1 vssd1 vccd1 vccd1 MuI._1217_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._4465__B MuI._0154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1305_ AuI._0490_ vssd1 vssd1 vccd1 vccd1 AuI._0503_ sky130_fd_sc_hd__inv_2
XFILLER_93_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0881__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3800__D MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5362_ MuI._2871_ MuI._0445_ vssd1 vssd1 vccd1 vccd1 MuI._1141_ sky130_fd_sc_hd__nand2_1
XAuI._1236_ AuI._0275_ AuI._0295_ AuI._0438_ vssd1 vssd1 vccd1 vccd1 AuI._0439_ sky130_fd_sc_hd__mux2_1
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4313_ MuI._3393_ MuI._3411_ MuI._3412_ vssd1 vssd1 vccd1 vccd1 MuI._3413_ sky130_fd_sc_hd__a21o_1
XFILLER_179_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07441__A _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5293_ MuI._0831_ MuI._1064_ vssd1 vssd1 vccd1 vccd1 MuI._1066_ sky130_fd_sc_hd__nor2_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _05708_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1167_ AuI._0274_ AuI._0293_ AuI._0373_ vssd1 vssd1 vccd1 vccd1 AuI._0374_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4244_ MuI._2704_ MuI._2803_ MuI._2539_ MuI._2495_ vssd1 vssd1 vccd1 vccd1 MuI._3344_
+ sky130_fd_sc_hd__and4_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5296__B MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1098_ AuI._0307_ AuI._0203_ AuI._0276_ vssd1 vssd1 vccd1 vccd1 AuI._0308_ sky130_fd_sc_hd__a21o_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4175_ MuI._3261_ MuI._3273_ MuI._3274_ vssd1 vssd1 vccd1 vccd1 MuI._3275_ sky130_fd_sc_hd__a21o_1
XANTENNA__11975__A2 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08840__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _00635_ _00636_ _00637_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__nand3_1
XANTENNA__13177__B2 _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09368__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12924__A1 _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3544__B MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _01878_ _01879_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a211o_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6816_ MuI._2710_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2739_ sky130_fd_sc_hd__and2b_1
XFILLER_115_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _01487_ _01488_ _01489_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__o21ba_1
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6747_ MuI._2659_ MuI._2664_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2665_ sky130_fd_sc_hd__mux2_1
XANTENNA__07616__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3959_ MuI._3055_ MuI._3058_ vssd1 vssd1 vccd1 vccd1 MuI._3059_ sky130_fd_sc_hd__xnor2_1
X_08853_ _01454_ _01469_ _01468_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a21o_1
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12241__B _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07804_ _02840_ _00421_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__nand2_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6678_ MuI._0787_ MuI._2582_ vssd1 vssd1 vccd1 vccd1 MuI._2589_ sky130_fd_sc_hd__nor2_1
XANTENNA__07335__B _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08784_ _01394_ _01401_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__xnor2_2
XFILLER_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5629_ MuI._1425_ MuI._1421_ MuI._1423_ vssd1 vssd1 vccd1 vccd1 MuI._1435_ sky130_fd_sc_hd__nor3_1
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07735_ _00350_ _00351_ _00352_ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__nand3_1
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI.pe._509_ AuI.pe._037_ AuI.pe._064_ AuI.pe._065_ AuI.pe._069_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[5\] sky130_fd_sc_hd__a31o_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._462__B AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07666_ _00280_ _00282_ _00283_ _06437_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__and4bb_1
XANTENNA_MuI._6243__A2 MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A2 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _02012_ _02014_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07351__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13072__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07597_ _06610_ _04918_ _00013_ _00010_ _00197_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__a32o_1
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09336_ _01835_ _01951_ _01950_ _01946_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a211o_1
XANTENNA__11304__C _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4006__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4006__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _06548_ _00035_ _04638_ _02291_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08292__B1 _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11601__A _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ _00820_ _00823_ _00821_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__o21ba_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _01690_ _01689_ _01688_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__o21ai_1
XFILLER_181_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11718__A2 _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08613__C _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08149_ _00764_ _00765_ _00750_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ _02550_ _05831_ _03802_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a31o_1
XFILLER_162_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4269__C MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _02784_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__nor2_1
X_11091_ _03306_ _02760_ _02722_ _02388_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10042_ _02020_ _06023_ _02075_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__nand3_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3470__A MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4493__A1 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input18_A a_operand[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09847__A1 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _04700_ _04810_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4493__B2 MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__B2 _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10944_ _02752_ _03506_ _03508_ _03682_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__a31o_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08357__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07261__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1021_ AuI._0147_ AuI._0232_ vssd1 vssd1 vccd1 vccd1 AuI._0233_ sky130_fd_sc_hd__nand2_2
X_10875_ _02712_ _03424_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__nand2_1
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11406__A1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ _05477_ _05479_ _05340_ _05344_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__o211ai_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6005__B MuI._1848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _00081_ _03082_ _00789_ _00086_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a22o_1
XFILLER_200_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08822__A2 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08092__A _00691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12476_ _05329_ _05330_ _05201_ _05219_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__a211o_1
XFILLER_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5980_ MuI._0775_ MuI._1820_ vssd1 vssd1 vccd1 vccd1 MuI._1821_ sky130_fd_sc_hd__and2_1
X_11427_ _03228_ _03282_ _00534_ _06525_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__and4_1
XFILLER_172_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10127__A _02801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4931_ MuI._0452_ MuI._0661_ MuI._0659_ vssd1 vssd1 vccd1 vccd1 MuI._0667_ sky130_fd_sc_hd__a21o_1
XAuI._0805_ net20 vssd1 vssd1 vccd1 vccd1 AuI._0025_ sky130_fd_sc_hd__inv_2
XANTENNA_MuI._6378__D MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ _03888_ _03892_ _04127_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__a211o_1
XANTENNA_AuI._0876__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._791_ AuI.pe._016_ AuI.pe._299_ vssd1 vssd1 vccd1 vccd1 AuI.pe._331_ sky130_fd_sc_hd__and2_1
XMuI._4862_ MuI.b_operand\[10\] MuI._2837_ MuI.a_operand\[10\] MuI.a_operand\[9\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0591_ sky130_fd_sc_hd__and4_1
X_10309_ _00703_ _00705_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__nor2_2
XFILLER_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _03979_ _03959_ _03961_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nand3_1
XANTENNA__12342__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6601_ MuI._2503_ vssd1 vssd1 vccd1 vccd1 MuI._2504_ sky130_fd_sc_hd__inv_2
XFILLER_112_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3813_ MuI._2911_ MuI._2912_ vssd1 vssd1 vccd1 vccd1 MuI._2913_ sky130_fd_sc_hd__xor2_2
XMuI._4793_ MuI._0386_ MuI._0388_ vssd1 vssd1 vccd1 vccd1 MuI._0516_ sky130_fd_sc_hd__xor2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13028_ _05918_ _05922_ _03133_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3744_ MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 MuI._2844_ sky130_fd_sc_hd__clkbuf_4
XMuI._6532_ MuI._1956_ MuI._2214_ MuI._2216_ MuI._2224_ vssd1 vssd1 vccd1 vccd1 MuI._2428_
+ sky130_fd_sc_hd__o31a_1
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07155__B _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6463_ MuI._2347_ MuI._2346_ vssd1 vssd1 vccd1 vccd1 MuI._2353_ sky130_fd_sc_hd__xor2_1
XMuI._3675_ MuI._1307_ MuI._2754_ MuI._2451_ MuI._2484_ vssd1 vssd1 vccd1 vccd1 MuI._2759_
+ sky130_fd_sc_hd__and4_1
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5414_ MuI._1192_ MuI._1193_ MuI._1198_ vssd1 vssd1 vccd1 vccd1 MuI._1199_ sky130_fd_sc_hd__a21o_1
XMuI._6394_ MuI._2100_ MuI._2270_ MuI._2269_ MuI._2276_ vssd1 vssd1 vccd1 vccd1 MuI._2277_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ _00135_ _00136_ _00137_ vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__and3_1
XANTENNA__09370__B _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5345_ MuI._1099_ MuI._1097_ MuI._1090_ vssd1 vssd1 vccd1 vccd1 MuI._1123_ sky130_fd_sc_hd__a21o_1
XFILLER_90_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07451_ _00044_ _00055_ _00068_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__a21o_1
XAuI._1219_ AuI._0330_ AuI._0222_ AuI._0234_ vssd1 vssd1 vccd1 vccd1 AuI._0423_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5276_ MuI._1044_ MuI._1045_ MuI._1036_ vssd1 vssd1 vccd1 vccd1 MuI._1047_ sky130_fd_sc_hd__a21o_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13398__B2 _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07382_ _06578_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__buf_4
XMuI._4227_ MuI._2671_ MuI._2975_ MuI._2976_ MuI._2616_ vssd1 vssd1 vccd1 vccd1 MuI._3327_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__08232__A1_N _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09121_ _06631_ _06630_ _04111_ _04176_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and4_1
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12517__A _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4158_ MuI._3161_ MuI._3164_ MuI._3163_ vssd1 vssd1 vccd1 vccd1 MuI._3258_ sky130_fd_sc_hd__o21ai_1
XFILLER_136_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09052_ _01586_ _01588_ _01668_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__and3_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08003_ _00620_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XMuI._4089_ MuI.b_operand\[7\] vssd1 vssd1 vccd1 vccd1 MuI._3189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08730__A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10384__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ _02340_ _02343_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__and2_1
XANTENNA__12252__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ _06630_ _00090_ _00093_ _06631_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22oi_1
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _02505_ _02506_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0928__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08836_ _01447_ _01448_ _01453_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__nand3_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08767_ _00029_ _04100_ _00271_ net120 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__a22o_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1410__A AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _00333_ _00332_ _00317_ _00298_ vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__o211a_1
XFILLER_199_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ _01311_ _01314_ _01277_ _01276_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__o211ai_1
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07081__A _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4227__A1 MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _00266_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4227__B2 MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07512__C _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _03338_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__xor2_2
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09452__A2_N _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _01928_ _01935_ _01936_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a21bo_1
XFILLER_210_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12061__A1 _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _02767_ _03302_ _02711_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12061__B2 _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ _05158_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__nor2_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3465__A MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ _05097_ _05098_ _05094_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__a21o_1
XFILLER_135_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09158__D net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _03967_ _03968_ _03969_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__a21o_1
XANTENNA__12364__A2 _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12192_ _04865_ _02728_ _02931_ FuI.Integer\[14\] vssd1 vssd1 vccd1 vccd1 _05026_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6152__A1 MuI._0482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _03893_ _03894_ _03721_ _03726_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__o211ai_1
XFILLER_123_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1570_ AuI._0701_ AuI._0742_ AuI._0746_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0747_
+ sky130_fd_sc_hd__o22a_1
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 ALU_Output[15] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 ALU_Output[25] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 ALU_Output[6] sky130_fd_sc_hd__buf_2
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11074_ _03819_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__xnor2_4
XANTENNA_MuI._4296__A MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0919__A1 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _00817_ _00818_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__and2_1
XFILLER_209_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11209__C _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6715__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3460_ MuI.b_operand\[24\] MuI.b_operand\[23\] MuI.b_operand\[26\] MuI.b_operand\[25\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0416_ sky130_fd_sc_hd__or4_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07703__B _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._520__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ net118 net117 _06461_ _05627_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__and4_1
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10927_ _03328_ _03662_ _03661_ _03296_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__a221o_1
XFILLER_72_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5130_ MuI._0859_ MuI._0860_ MuI._0861_ vssd1 vssd1 vccd1 vccd1 MuI._0886_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1004_ net40 net8 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0216_ sky130_fd_sc_hd__mux2_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10858_ _03571_ _03573_ _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a21oi_2
XFILLER_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5061_ MuI._0168_ MuI._3371_ MuI._0808_ MuI._0809_ vssd1 vssd1 vccd1 vccd1 MuI._0810_
+ sky130_fd_sc_hd__and4_1
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4012_ MuI.b_operand\[21\] MuI._2791_ MuI._2787_ MuI.b_operand\[22\] vssd1 vssd1
+ vccd1 vccd1 MuI._3112_ sky130_fd_sc_hd__a22o_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _03380_ _03412_ _03413_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__and3_1
XFILLER_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ _02613_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__xor2_2
XFILLER_185_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09349__C _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08008__B1 _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12459_ net113 _03432_ _06489_ _05498_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__and4_1
XFILLER_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5963_ MuI._0769_ MuI._1800_ MuI._1788_ MuI._1787_ vssd1 vssd1 vccd1 vccd1 MuI._1803_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_160_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11563__B1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4914_ MuI._0607_ MuI._0609_ MuI._0648_ MuI._0455_ vssd1 vssd1 vccd1 vccd1 MuI._0649_
+ sky130_fd_sc_hd__a211o_1
XFILLER_113_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13168__A _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5894_ MuI._1164_ MuI._0246_ MuI._0420_ MuI._0746_ vssd1 vssd1 vccd1 vccd1 MuI._1727_
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09365__B _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12072__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4845_ MuI._0560_ MuI._0569_ MuI._0571_ vssd1 vssd1 vccd1 vccd1 MuI._0573_ sky130_fd_sc_hd__or3_1
XANTENNA__07166__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _04896_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._3901__B1 MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12222__D _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4776_ MuI._0456_ MuI._0495_ MuI._0496_ vssd1 vssd1 vccd1 vccd1 MuI._0497_ sky130_fd_sc_hd__a21bo_1
X_09670_ _02256_ _02308_ _02304_ _02307_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__o211a_1
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06882_ net125 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__clkbuf_4
XMuI._6515_ MuI._2408_ MuI._2400_ vssd1 vssd1 vccd1 vccd1 MuI._2410_ sky130_fd_sc_hd__and2b_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3727_ MuI._2826_ MuI._0603_ MuI._2385_ MuI._2330_ vssd1 vssd1 vccd1 vccd1 MuI._2827_
+ sky130_fd_sc_hd__and4_1
XFILLER_95_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08621_ _01084_ _01238_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3658_ MuI._2528_ vssd1 vssd1 vccd1 vccd1 MuI._2594_ sky130_fd_sc_hd__buf_2
XMuI._6446_ MuI._2295_ MuI._2329_ MuI._2320_ MuI._2328_ vssd1 vssd1 vccd1 vccd1 MuI._2334_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_208_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08552_ _01150_ _01169_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__or2_1
X_07503_ _00107_ _00108_ _00120_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__a21oi_4
XANTENNA_MuI._4209__A1 MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6377_ MuI._0603_ MuI._2594_ MuI._2797_ MuI._2826_ vssd1 vssd1 vccd1 vccd1 MuI._2258_
+ sky130_fd_sc_hd__a22oi_1
XMuI._3589_ MuI._1813_ MuI._0515_ MuI._1329_ vssd1 vssd1 vccd1 vccd1 MuI._1835_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4209__B2 MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07332__C _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _01099_ _01100_ _03163_ _00303_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__and4bb_1
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5328_ MuI._1101_ MuI._1102_ MuI._1103_ vssd1 vssd1 vccd1 vccd1 MuI._1104_ sky130_fd_sc_hd__nand3_1
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07434_ _00045_ _00051_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__or2_1
XFILLER_51_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3968__B1 MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4091__D MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5765__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5259_ MuI._1024_ MuI._1025_ MuI._1026_ vssd1 vssd1 vccd1 vccd1 MuI._1028_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12043__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07365_ _05434_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__buf_4
XFILLER_176_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12247__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _01418_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__nor2_2
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07296_ _06588_ _06595_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _01203_ _01652_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__or2_1
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3716__C MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09275__B _01891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07076__A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09937_ _02336_ _02337_ _02325_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__o21a_1
XANTENNA_AuI.pe._735__C1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__A1 _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__D _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09868_ _02479_ _02492_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07226__D net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _01415_ _01436_ _01410_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07804__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13059__B1 _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _02441_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__nor2b_1
XANTENNA_MuI._4786__A2_N MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _04634_ _02892_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._4999__A2 MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5659__B MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4563__B MuI._0208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__D net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07289__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__xor2_4
XFILLER_26_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _03429_ _03430_ _03431_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nand3_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _04359_ _04487_ _04488_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08635__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _05853_ _02745_ _02722_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__a21o_1
X_10643_ _02980_ _00036_ _04649_ _02983_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a22o_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12585__A2 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ _06245_ _06244_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__nor2_1
XFILLER_182_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _03137_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10596__A1 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__C _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _05154_ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__and2_1
XFILLER_182_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _06200_ _06201_ _06199_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a21o_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12244_ _05081_ _05082_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__xnor2_4
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08370__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11545__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1622_ AuI.pe.Significand\[18\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0790_
+ sky130_fd_sc_hd__or2_1
X_12175_ _02447_ _05008_ _02581_ _04881_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a211o_1
XFILLER_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08410__B1 _01026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__A1 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11126_ _00502_ _04380_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__nand2_1
XFILLER_123_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1553_ AuI._0732_ AuI._0648_ vssd1 vssd1 vccd1 vccd1 AuI._0733_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4630_ MuI._0334_ MuI._0332_ vssd1 vssd1 vccd1 vccd1 MuI._0336_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1014__A0 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11848__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _02539_ _03257_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__nand2_1
XAuI._1484_ AuI._0524_ AuI._0527_ vssd1 vssd1 vccd1 vccd1 AuI._0670_ sky130_fd_sc_hd__and2_1
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11848__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4561_ MuI._0258_ MuI._0259_ vssd1 vssd1 vccd1 vccd1 MuI._0260_ sky130_fd_sc_hd__nor2_1
XAuI.pe._490_ AuI.pe._037_ AuI.pe._047_ AuI.pe._049_ AuI.pe._052_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[3\] sky130_fd_sc_hd__a31o_1
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07516__A2 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _02671_ _02674_ _02675_ _02662_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__o211a_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__C _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6300_ MuI._0878_ MuI._1494_ MuI._2172_ vssd1 vssd1 vccd1 vccd1 MuI._2173_ sky130_fd_sc_hd__and3_1
XMuI._3512_ MuI._0724_ MuI._0977_ vssd1 vssd1 vccd1 vccd1 MuI._0988_ sky130_fd_sc_hd__or2_1
XMuI._4492_ MuI._2850_ MuI._2495_ vssd1 vssd1 vccd1 vccd1 MuI._0184_ sky130_fd_sc_hd__nand2_1
XANTENNA__10140__A _02815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6231_ MuI._2095_ MuI._2096_ vssd1 vssd1 vccd1 vccd1 MuI._2097_ sky130_fd_sc_hd__xnor2_1
XMuI._3443_ MuI.a_operand\[26\] MuI.b_operand\[26\] vssd1 vssd1 vccd1 vccd1 MuI._0229_
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11959_ _04772_ _04773_ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nand3b_1
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6162_ MuI._1021_ MuI._2550_ MuI._2517_ MuI._0779_ vssd1 vssd1 vccd1 vccd1 MuI._2021_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12993__C _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5939__A1 MuI._0725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5113_ MuI._2765_ MuI.a_operand\[9\] MuI._3306_ MuI._3307_ vssd1 vssd1 vccd1
+ vccd1 MuI._0868_ sky130_fd_sc_hd__and4_1
XMuI._6093_ MuI._1943_ MuI._1944_ vssd1 vssd1 vccd1 vccd1 MuI._1946_ sky130_fd_sc_hd__nor2_1
XFILLER_193_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5044_ MuI._3303_ MuI._0791_ MuI._3302_ vssd1 vssd1 vccd1 vccd1 MuI._0792_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ _03733_ _03906_ _06449_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _04607_ _06284_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and2_1
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10339__A1 _00734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5946_ MuI._1740_ MuI._1751_ vssd1 vssd1 vccd1 vccd1 MuI._1784_ sky130_fd_sc_hd__or2_1
Xfanout106 net67 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_6
XAuI.pe._826_ AuI.operand_a\[27\] AuI.pe._273_ AuI.pe._360_ AuI.pe._362_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._363_ sky130_fd_sc_hd__a22o_1
Xfanout117 net47 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_4
XANTENNA__08952__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5877_ MuI._1705_ MuI._1706_ MuI._1631_ MuI._1650_ vssd1 vssd1 vccd1 vccd1 MuI._1708_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_102_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout128 net26 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_4
X_07983_ _00313_ _00314_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__B _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._757_ AuI.pe._158_ AuI.pe._391_ AuI.pe._118_ AuI.pe.significand\[12\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._301_ sky130_fd_sc_hd__a22o_1
XMuI._4828_ MuI.a_operand\[17\] MuI.b_operand\[1\] MuI._0018_ MuI.a_operand\[18\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0554_ sky130_fd_sc_hd__a22oi_1
X_09722_ _06545_ _04046_ _02352_ _02351_ _02350_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a32o_1
XANTENNA__11839__A1 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ _04714_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__buf_4
XANTENNA__11839__B2 _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._688_ AuI.pe._125_ AuI.pe._097_ AuI.pe._233_ AuI.pe._235_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._236_ sky130_fd_sc_hd__a211o_1
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4086__D MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4759_ MuI.b_operand\[10\] MuI._2837_ MuI._0477_ MuI.a_operand\[10\] vssd1 vssd1
+ vccd1 vccd1 MuI._0478_ sky130_fd_sc_hd__and4_1
X_09653_ _02273_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__nor2_1
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06865_ _03971_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__buf_4
XFILLER_110_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11146__A _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _06479_ _06480_ _06581_ _05101_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__and4_1
XANTENNA__07343__B net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09584_ _02166_ _02218_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10050__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06796_ _03228_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1308__A1 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6429_ MuI._1939_ MuI._2311_ MuI._2313_ MuI._2314_ vssd1 vssd1 vccd1 vccd1 MuI._2315_
+ sky130_fd_sc_hd__a211oi_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _01142_ _01151_ _01152_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__a21o_1
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08466_ net121 _04445_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__nand2_1
XFILLER_211_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ net6 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__buf_4
XANTENNA__12016__A1 _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _01007_ _01008_ _01014_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__a21oi_2
XFILLER_211_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3727__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _06646_ _06647_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nand3_1
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ net133 vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12705__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ _01539_ _01543_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__or2b_1
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10290_ _00729_ _00732_ _00730_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__o21bai_1
XFILLER_145_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3743__A MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__C1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07534__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12931_ _05817_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__xnor2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08349__B _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _05661_ _05663_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__o21ai_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11813_ _04614_ _04617_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__nor2_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12793_ _02854_ _05582_ _02868_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__a21o_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09120__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09120__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11744_ _04525_ _04526_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a21o_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ _04428_ _04429_ _04469_ _04470_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__o211ai_4
XANTENNA__08084__B _00698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _06289_ _06292_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__o21a_1
X_10626_ _03744_ _04197_ _03149_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nand3_1
XFILLER_186_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__A2 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5149__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13345_ _06254_ _06255_ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__o21a_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _03256_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__xnor2_2
XAuI._0984_ AuI._0115_ AuI._0194_ AuI._0195_ AuI._0148_ vssd1 vssd1 vccd1 vccd1 AuI._0196_
+ sky130_fd_sc_hd__or4_1
XFILLER_170_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _06102_ _06184_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__or2_1
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10488_ _03189_ _03190_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a21o_1
XMuI._5800_ MuI._1620_ MuI._1621_ MuI._1608_ vssd1 vssd1 vccd1 vccd1 MuI._1623_ sky130_fd_sc_hd__a21o_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09187__A1 _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3653__A MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6780_ MuI._2588_ MuI._2597_ MuI._2601_ vssd1 vssd1 vccd1 vccd1 MuI._2701_ sky130_fd_sc_hd__a21oi_1
X_12227_ _04925_ _04927_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nand2_1
XMuI._3992_ MuI._3091_ MuI._2860_ MuI._3050_ MuI._3049_ vssd1 vssd1 vccd1 vccd1 MuI._3092_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10135__A _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5731_ MuI._1478_ MuI._1545_ MuI._1546_ vssd1 vssd1 vccd1 vccd1 MuI._1547_ sky130_fd_sc_hd__nand3_1
XFILLER_151_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1605_ AuI._0673_ AuI._0775_ vssd1 vssd1 vccd1 vccd1 AuI._0776_ sky130_fd_sc_hd__nand2_1
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12730__A2 _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12158_ _04987_ _04988_ _04853_ _04905_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__o211a_1
XAuI.pe._611_ AuI.pe._380_ AuI.pe._149_ AuI.pe._395_ vssd1 vssd1 vccd1 vccd1 AuI.pe._164_
+ sky130_fd_sc_hd__and3_2
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0884__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5662_ MuI._1467_ MuI._1470_ vssd1 vssd1 vccd1 vccd1 MuI._1471_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11109_ _03591_ _03594_ _03734_ _03735_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__o211a_1
XFILLER_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1536_ AuI._0702_ vssd1 vssd1 vccd1 vccd1 AuI._0719_ sky130_fd_sc_hd__buf_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3868__C1 MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _04913_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._542_ AuI.pe._055_ AuI.pe._079_ AuI.pe._097_ AuI.pe._020_ AuI.pe._099_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._100_ sky130_fd_sc_hd__a221o_1
XFILLER_65_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4613_ MuI.b_operand\[21\] MuI._0111_ MuI._0315_ MuI._2826_ vssd1 vssd1 vccd1
+ vccd1 MuI._0318_ sky130_fd_sc_hd__a22o_1
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07444__A _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5593_ MuI._1379_ MuI._1380_ vssd1 vssd1 vccd1 vccd1 MuI._1396_ sky130_fd_sc_hd__nor2_1
XAuI._1467_ AuI._0320_ AuI._0323_ vssd1 vssd1 vccd1 vccd1 AuI._0653_ sky130_fd_sc_hd__or2_1
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._473_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._037_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4544_ MuI._2826_ MuI._0603_ MuI._3372_ MuI._0112_ vssd1 vssd1 vccd1 vccd1 MuI._0242_
+ sky130_fd_sc_hd__and4_1
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1398_ AuI._0258_ AuI._0584_ AuI._0585_ AuI._0586_ vssd1 vssd1 vccd1 vccd1 AuI._0588_
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4475_ MuI._0165_ MuI._0033_ vssd1 vssd1 vccd1 vccd1 MuI._0166_ sky130_fd_sc_hd__xnor2_2
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6214_ MuI._1971_ MuI._1973_ MuI._1972_ vssd1 vssd1 vccd1 vccd1 MuI._2079_ sky130_fd_sc_hd__o21bai_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3426_ MuI.a_operand\[24\] MuI.a_operand\[26\] MuI.a_operand\[25\] vssd1 vssd1
+ vccd1 vccd1 MuI._0043_ sky130_fd_sc_hd__and3_1
X_08320_ _00614_ _00616_ _00617_ _00615_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a22o_1
XANTENNA__10114__A_N _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6145_ MuI._1999_ MuI._1998_ vssd1 vssd1 vccd1 vccd1 MuI._2003_ sky130_fd_sc_hd__and2b_1
X_08251_ _00866_ _00867_ _00857_ _00862_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__a211o_1
XANTENNA__07673__A1 _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07673__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__B1 _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ net110 vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__buf_4
XMuI._6076_ MuI._1852_ MuI._1858_ vssd1 vssd1 vccd1 vccd1 MuI._1927_ sky130_fd_sc_hd__or2b_1
XANTENNA__11132__C _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _00798_ _00799_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._5465__D MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5027_ MuI._0709_ MuI._0737_ MuI._0739_ vssd1 vssd1 vccd1 vccd1 MuI._0773_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI.pe._650__A1 AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._650__B2 AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07133_ net112 vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__buf_2
XFILLER_118_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout118_A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07064_ _04068_ _06067_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__and2_1
XFILLER_133_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07619__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07728__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5929_ MuI._1761_ MuI._1764_ vssd1 vssd1 vccd1 vccd1 MuI._1765_ sky130_fd_sc_hd__or2_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._809_ AuI.pe._346_ AuI.pe._336_ AuI.pe._347_ vssd1 vssd1 vccd1 vccd1 AuI.pe._348_
+ sky130_fd_sc_hd__or3_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _00580_ _00581_ _00583_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__or3_1
XFILLER_56_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__B _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09705_ _02301_ _02300_ _02293_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a21o_1
X_06917_ _04531_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__clkbuf_4
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4394__A MuI._0075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07897_ _00504_ _06450_ _00514_ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__o21a_1
X_09636_ _02231_ _02230_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__nor2_1
XANTENNA__11693__C1 _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1607__B1_N AuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ net61 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__clkbuf_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4544__D MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _02197_ _02198_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__o21bai_1
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06779_ net118 vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__buf_4
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08518_ _01134_ _01133_ _01119_ _01066_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__o211a_1
XFILLER_196_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ _02111_ _02116_ _02110_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a21bo_1
XFILLER_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3738__A MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07664__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08449_ _01065_ _01064_ _01050_ _01017_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__a211o_1
XANTENNA__07664__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFuI._153_ FuI.a_operand\[23\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[23\] sky130_fd_sc_hd__clkbuf_1
XFILLER_184_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _04230_ _04231_ _04236_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__o21bai_1
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._084_ FuI._038_ FuI._044_ FuI._039_ vssd1 vssd1 vccd1 vccd1 FuI._048_ sky130_fd_sc_hd__and3_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ _00805_ _00804_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__and2b_1
XANTENNA__07416__A1 _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ _04162_ _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07416__B2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08632__B _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _03809_ _05595_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nand3_1
X_10342_ _03033_ _03034_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__and2b_1
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _03669_ _05660_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__nand2_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07248__B _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ _03733_ _04068_ _00684_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__nand3_1
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _03217_ _03271_ _06562_ _06476_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__and4_1
XANTENNA__12712__A2 _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A b_operand[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1321_ AuI._0503_ AuI._0504_ AuI._0515_ AuI._0486_ vssd1 vssd1 vccd1 vccd1 AuI._0518_
+ sky130_fd_sc_hd__or4b_2
XANTENNA__07264__A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08079__B _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12914_ _05708_ _05709_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__a21oi_1
XAuI._1252_ net6 net38 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0454_ sky130_fd_sc_hd__mux2_2
XFILLER_207_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5067__A1 MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5067__B2 MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07352__B1 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12845_ _05726_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__nor2_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1183_ AuI._0153_ vssd1 vssd1 vccd1 vccd1 AuI._0389_ sky130_fd_sc_hd__buf_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4260_ MuI._3239_ MuI._3359_ vssd1 vssd1 vccd1 vccd1 MuI._3360_ sky130_fd_sc_hd__nor2_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _05651_ _05652_ _05610_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o21ai_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4191_ MuI._2825_ MuI._2831_ MuI._2827_ vssd1 vssd1 vccd1 vccd1 MuI._3291_ sky130_fd_sc_hd__o21ba_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3648__A MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ _04522_ _04523_ _04524_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a21o_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _00345_ _04918_ _04450_ _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a22o_1
XANTENNA_AuI._0879__A net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ _02714_ _02881_ _03320_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a21o_1
XANTENNA__11203__A2 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12400__B2 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ _06608_ _03449_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13328_ _06237_ _06238_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__or2_1
XFILLER_171_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09357__C net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0967_ net47 net15 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0179_ sky130_fd_sc_hd__mux2_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6832_ MuI._2747_ vssd1 vssd1 vccd1 vccd1 MuI.result\[8\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08261__C _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07158__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ _02827_ _02875_ _06108_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__or3_1
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0898_ net128 net58 vssd1 vssd1 vccd1 vccd1 AuI._0118_ sky130_fd_sc_hd__or2b_1
XANTENNA__12999__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__B1 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6763_ MuI._2681_ vssd1 vssd1 vccd1 vccd1 MuI._2683_ sky130_fd_sc_hd__dlymetal6s2s_1
XMuI._3975_ MuI._3072_ MuI._3073_ MuI._3074_ vssd1 vssd1 vccd1 vccd1 MuI._3075_ sky130_fd_sc_hd__and3_1
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5714_ MuI._2605_ MuI._3262_ MuI._0020_ MuI._2852_ vssd1 vssd1 vccd1 vccd1 MuI._1529_
+ sky130_fd_sc_hd__a22oi_2
X_07820_ _00186_ _00372_ _00436_ _00437_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__o211ai_1
XMuI._6694_ MuI._1996_ MuI._2606_ vssd1 vssd1 vccd1 vccd1 MuI._2607_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6810__B_N MuI._2733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__D net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5645_ MuI._1294_ MuI._1331_ MuI._1332_ MuI._1371_ vssd1 vssd1 vccd1 vccd1 MuI._1453_
+ sky130_fd_sc_hd__and4_1
XANTENNA_AuI.pe._699__B2 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1519_ AuI._0656_ AuI._0653_ vssd1 vssd1 vccd1 vccd1 AuI._0704_ sky130_fd_sc_hd__or2b_1
X_07751_ _00366_ _00367_ _00334_ _00339_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__o211ai_2
XAuI.pe._525_ AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 AuI.pe._084_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4645__C MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _02216_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__and3_1
XMuI._5576_ MuI._1356_ MuI._1347_ MuI._1355_ vssd1 vssd1 vccd1 vccd1 MuI._1377_ sky130_fd_sc_hd__nand3_1
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07682_ _00299_ _00231_ _00287_ _00267_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__and4_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._456_ AuI.pe._021_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4527_ MuI._0220_ MuI._0222_ vssd1 vssd1 vccd1 vccd1 MuI._0223_ sky130_fd_sc_hd__nand2_1
X_09421_ _01847_ _01881_ _02040_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__and3_1
XANTENNA__11400__B_N _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4458_ MuI._0145_ MuI._0146_ vssd1 vssd1 vccd1 vccd1 MuI._0147_ sky130_fd_sc_hd__or2_1
X_09352_ _01968_ _01969_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07621__B _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5757__B MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ _00237_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__buf_6
XFILLER_61_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3558__A MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4389_ MuI._0069_ MuI._0070_ MuI._0059_ MuI._0063_ vssd1 vssd1 vccd1 vccd1 MuI._0072_
+ sky130_fd_sc_hd__o211ai_1
X_09283_ _01899_ _01900_ _02712_ _04111_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__and4bb_1
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6128_ MuI._1981_ MuI._1983_ vssd1 vssd1 vccd1 vccd1 MuI._1984_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08234_ _06578_ _02647_ _06602_ _06604_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__and4_1
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6059_ MuI._1849_ MuI._1907_ vssd1 vssd1 vccd1 vccd1 MuI._1908_ sky130_fd_sc_hd__xnor2_2
XFILLER_193_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ net128 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07116_ _05724_ _06414_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__and2_1
XANTENNA__07949__A2 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08096_ _00422_ _00424_ _00425_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__o21bai_1
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07047_ _05928_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[30\] sky130_fd_sc_hd__clkbuf_2
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1531__B1_N AuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09564__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5297__A1 MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _01508_ _01509_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__or4bb_1
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _02840_ _00059_ _00565_ _00566_ _00555_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a32o_2
XANTENNA__12458__B2 _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5049__A1 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ _00678_ _00085_ _00047_ _03539_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__a22o_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5049__B2 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__D net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _02253_ _02254_ _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__nor3_2
XFILLER_189_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10891_ _03622_ _03623_ _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand3b_1
XFILLER_204_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _01206_ _03444_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nand2_1
XFILLER_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11969__B1 _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3468__A MuI._0482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _05297_ _05296_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or2b_1
XFILLER_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _04291_ _04292_ _04253_ _04254_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__a211o_1
XFILLER_211_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _05130_ _05131_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__xor2_1
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._136_ FuI._020_ net142 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[7\] sky130_fd_sc_hd__dlxtn_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11443_ _04045_ _04048_ _04218_ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__a211oi_1
XFILLER_184_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09458__B _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08362__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._067_ FuI.a_operand\[27\] net105 FuI._033_ FuI._034_ vssd1 vssd1 vccd1 vccd1
+ FuI._035_ sky130_fd_sc_hd__a31o_1
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07259__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0821_ AuI._0038_ net15 vssd1 vssd1 vccd1 vccd1 AuI._0041_ sky130_fd_sc_hd__or2_1
X_11374_ _04145_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__nor2_2
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10944__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _02841_ _06012_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__or2_1
XFILLER_153_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10325_ _03014_ _03015_ _03007_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__a21o_1
XFILLER_152_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6010__C MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09474__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _05877_ _05879_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and2b_1
X_10256_ _04004_ _02941_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nor2_1
XFILLER_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3760_ MuI._2796_ vssd1 vssd1 vccd1 vccd1 MuI._2860_ sky130_fd_sc_hd__clkbuf_4
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _02866_ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__nor2_2
XANTENNA__10178__B_N _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3650__B MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3691_ MuI._2790_ vssd1 vssd1 vccd1 vccd1 MuI._2791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6019__A MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5430_ MuI._1139_ MuI._1151_ MuI._1150_ vssd1 vssd1 vccd1 vccd1 MuI._1216_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09314__A1 _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__B2 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1304_ AuI._0486_ AuI._0490_ AuI._0501_ vssd1 vssd1 vccd1 vccd1 AuI._0502_ sky130_fd_sc_hd__a21o_1
XFILLER_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0881__B net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5361_ MuI._1125_ MuI._1127_ MuI._1124_ vssd1 vssd1 vccd1 vccd1 MuI._1140_ sky130_fd_sc_hd__o21ba_1
XFILLER_90_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1235_ AuI._0263_ vssd1 vssd1 vccd1 vccd1 AuI._0438_ sky130_fd_sc_hd__clkbuf_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4312_ MuI._3410_ MuI._3408_ vssd1 vssd1 vccd1 vccd1 MuI._3412_ sky130_fd_sc_hd__and2b_1
XFILLER_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5292_ MuI._2851_ MuI._0320_ MuI._0829_ MuI._0830_ vssd1 vssd1 vccd1 vccd1 MuI._1064_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_179_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12828_ _05620_ _05622_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nand2_1
XAuI._1166_ AuI._0176_ AuI._0236_ AuI._0198_ AuI._0307_ vssd1 vssd1 vccd1 vccd1 AuI._0373_
+ sky130_fd_sc_hd__a31o_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4243_ MuI._2919_ MuI._2539_ MuI._2789_ MuI._2800_ vssd1 vssd1 vccd1 vccd1 MuI._3343_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08825__B1 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _05633_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__xnor2_1
XAuI._1097_ AuI._0223_ vssd1 vssd1 vccd1 vccd1 AuI._0307_ sky130_fd_sc_hd__buf_2
XMuI._4174_ MuI._3270_ MuI._3272_ vssd1 vssd1 vccd1 vccd1 MuI._3274_ sky130_fd_sc_hd__and2_1
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11898__B _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09368__B _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4971__B1 MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12924__A2 _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07169__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6712__A1 MuI._2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09970_ _01848_ _01849_ _01878_ _01879_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__o211ai_2
XFILLER_115_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0947__B_N AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6815_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2738_ sky130_fd_sc_hd__clkbuf_2
XFILLER_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08921_ _01499_ _01501_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__nor2_1
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06801__A _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6746_ MuI._2662_ MuI._2663_ vssd1 vssd1 vccd1 vccd1 MuI._2664_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08356__A2 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3958_ MuI._3056_ MuI._3057_ vssd1 vssd1 vccd1 vccd1 MuI._3058_ sky130_fd_sc_hd__xor2_1
X_08852_ _01454_ _01468_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nand3_2
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07616__B _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12241__C _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07803_ _06584_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__buf_4
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6677_ MuI._2577_ MuI._2580_ MuI._2587_ vssd1 vssd1 vccd1 vccd1 MuI._2588_ sky130_fd_sc_hd__and3_1
XMuI._3889_ MuI._2981_ MuI._2982_ MuI._2987_ vssd1 vssd1 vccd1 vccd1 MuI._2989_ sky130_fd_sc_hd__a21o_1
X_08783_ _01395_ _01400_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5628_ MuI._1431_ MuI._1427_ vssd1 vssd1 vccd1 vccd1 MuI._1434_ sky130_fd_sc_hd__xor2_1
XFILLER_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07734_ _00348_ _00349_ _00344_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a21o_1
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._541__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI.pe._508_ AuI.pe._020_ AuI.pe._066_ AuI.pe._054_ AuI.pe._029_ AuI.pe._068_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._069_ sky130_fd_sc_hd__a221o_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5559_ MuI._1344_ MuI._1345_ MuI._1357_ vssd1 vssd1 vccd1 vccd1 MuI._1358_ sky130_fd_sc_hd__a21oi_1
X_07665_ net55 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__buf_4
XFILLER_198_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12860__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._439_ AuI.pe.significand\[22\] AuI.pe._005_ vssd1 vssd1 vccd1 vccd1 AuI.pe._006_
+ sky130_fd_sc_hd__and2_1
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _01921_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__nand2_1
XANTENNA__11154__A _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07351__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07596_ _00109_ _00112_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__or2b_1
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _01921_ _01922_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__xor2_1
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12612__A1 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__D _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _01776_ _01778_ _01777_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08292__A1 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4006__A2 MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08292__B2 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08217_ _00819_ _00833_ _00834_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__nand3_4
XANTENNA__11601__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09197_ _01690_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__or3_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08148_ _00750_ _00764_ _00765_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__and3_1
XANTENNA__08613__D _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _00283_ _00259_ _00694_ _00695_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__nand4_2
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10110_ _04467_ _02550_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__and2b_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07807__A _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4269__D MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11090_ _02760_ _03838_ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__o21a_1
XFILLER_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3751__A MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _02710_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__buf_2
XANTENNA__11329__A _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._532__B1 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11992_ _04768_ _04769_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a22o_1
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4493__A2 MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09847__A2 _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07542__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ _03134_ _03666_ _03667_ _03670_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__a311o_1
XFILLER_44_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1020_ AuI._0207_ AuI._0100_ vssd1 vssd1 vccd1 vccd1 AuI._0232_ sky130_fd_sc_hd__or2b_1
X_10874_ _06585_ _06583_ _05638_ _06537_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__and4_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12613_ _05340_ _05344_ _05477_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__a211oi_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0921__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__B1 _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12544_ _05403_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xnor2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12475_ _05201_ _05219_ _05329_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o211ai_4
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._119_ FuI._038_ FuI._024_ vssd1 vssd1 vccd1 vccd1 FuI._030_ sky130_fd_sc_hd__nand2_1
XFILLER_126_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _00727_ _00423_ _05198_ _00728_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a22oi_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10127__B _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4930_ MuI._0664_ MuI._0665_ vssd1 vssd1 vccd1 vccd1 MuI._0666_ sky130_fd_sc_hd__or2b_1
XFILLER_126_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11357_ _04125_ _04126_ _04115_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._790_ AuI.pe._318_ AuI.pe._327_ AuI.pe._326_ vssd1 vssd1 vccd1 vccd1 AuI.pe._330_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_180_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4861_ MuI._0587_ MuI._0586_ MuI._0585_ MuI._0572_ vssd1 vssd1 vccd1 vccd1 MuI._0590_
+ sky130_fd_sc_hd__o211a_1
X_10308_ _02996_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__nor2_1
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11288_ _04050_ _04051_ _03943_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a21oi_1
XMuI._6600_ MuI._0141_ MuI._2502_ vssd1 vssd1 vccd1 vccd1 MuI._2503_ sky130_fd_sc_hd__xor2_2
XANTENNA__12342__B _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3812_ MuI._2839_ MuI._2847_ vssd1 vssd1 vccd1 vccd1 MuI._2912_ sky130_fd_sc_hd__or2b_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3661__A MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13027_ _05918_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__nand2_1
XMuI._4792_ MuI._0511_ MuI._0513_ vssd1 vssd1 vccd1 vccd1 MuI._0514_ sky130_fd_sc_hd__and2_1
X_10239_ _03842_ _02875_ _02826_ _02915_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__o221ai_4
XFILLER_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10143__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4476__B MuI._0166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6531_ MuI._2411_ MuI._2413_ vssd1 vssd1 vccd1 vccd1 MuI._2427_ sky130_fd_sc_hd__and2_1
XMuI._3743_ MuI._2055_ vssd1 vssd1 vccd1 vccd1 MuI._2843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0892__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07155__C _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6462_ MuI._2326_ MuI._2350_ vssd1 vssd1 vccd1 vccd1 MuI._2351_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3674_ MuI.b_operand\[15\] vssd1 vssd1 vccd1 vccd1 MuI._2754_ sky130_fd_sc_hd__buf_2
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5413_ MuI._1194_ MuI._1195_ MuI._1196_ vssd1 vssd1 vccd1 vccd1 MuI._1198_ sky130_fd_sc_hd__o21bai_1
XFILLER_35_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6393_ MuI._2271_ MuI._1975_ MuI._2272_ vssd1 vssd1 vccd1 vccd1 MuI._2276_ sky130_fd_sc_hd__a21oi_2
XFILLER_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3692__B1 MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4492__A MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5344_ MuI._1099_ MuI._1090_ MuI._1097_ vssd1 vssd1 vccd1 vccd1 MuI._1122_ sky130_fd_sc_hd__nand3_1
X_07450_ _00056_ _00067_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__xnor2_1
XAuI._1218_ AuI._0421_ vssd1 vssd1 vccd1 vccd1 AuI._0422_ sky130_fd_sc_hd__clkbuf_2
XFILLER_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._826__A1 AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5275_ MuI._1036_ MuI._1044_ MuI._1045_ vssd1 vssd1 vccd1 vccd1 MuI._1046_ sky130_fd_sc_hd__nand3_1
XANTENNA__13398__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5100__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07381_ _06579_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__buf_4
XAuI._1149_ AuI._0262_ AuI._0330_ AuI._0356_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0357_
+ sky130_fd_sc_hd__o31a_1
XFILLER_188_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4226_ MuI._2528_ MuI._2850_ vssd1 vssd1 vccd1 vccd1 MuI._3326_ sky130_fd_sc_hd__nand2_1
X_09120_ _00011_ _04111_ _00272_ _06631_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._3995__B2 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4157_ MuI._3256_ MuI._3210_ vssd1 vssd1 vccd1 vccd1 MuI._3257_ sky130_fd_sc_hd__xnor2_2
XFILLER_176_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _01586_ _01588_ _01668_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08002_ _00614_ _00618_ _00588_ _00619_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__a211o_1
XFILLER_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4088_ MuI._2878_ MuI._3183_ MuI._3187_ vssd1 vssd1 vccd1 vccd1 MuI._3188_ sky130_fd_sc_hd__a21o_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08730__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A2 _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _02614_ _02616_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__and2_1
XANTENNA__13348__B _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _02754_ _02797_ _04358_ _00083_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__and4_1
X_09884_ _02302_ _03917_ _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__and3_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6729_ MuI._2459_ MuI._2644_ vssd1 vssd1 vccd1 vccd1 MuI._2645_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._754__A AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _01449_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ net120 net44 _04100_ _04165_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__and4_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07362__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _00298_ _00317_ _00332_ _00333_ vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__a211oi_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _01276_ _01277_ _01314_ _01311_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__a211o_1
XANTENNA__10500__B _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ net124 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4227__A2 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07512__D _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._817__A1 AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07579_ _04961_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__buf_4
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _01929_ _01934_ _01930_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__nand3_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10590_ _02559_ _02753_ _02532_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__o21a_1
XANTENNA__12061__A2 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06706__A _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _01865_ _01864_ _01851_ _01644_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a211oi_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0864__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _05094_ _05097_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nand3_2
XFILLER_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ _03967_ _03968_ _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__nand3_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11021__B1 _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _04800_ _04642_ _05022_ _05023_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a211o_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ _03721_ _03726_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._6152__A2 MuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09455__C _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 ALU_Output[16] sky130_fd_sc_hd__buf_2
XANTENNA_MuI._3481__A MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 ALU_Output[26] sky130_fd_sc_hd__buf_2
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11073_ _03558_ _03646_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 ALU_Output[7] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10024_ _02679_ _02683_ _02693_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__and3_1
XANTENNA_input30_A a_operand[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5112__B1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11209__D _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07272__A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11088__B1 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11975_ _00462_ _05563_ _05638_ _00237_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a22oi_2
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ _03331_ _03484_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_17_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1003_ AuI._0190_ AuI._0191_ AuI._0214_ vssd1 vssd1 vccd1 vccd1 AuI._0215_ sky130_fd_sc_hd__or3b_1
XFILLER_189_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10857_ _03578_ _03587_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._6731__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5060_ MuI._2868_ MuI.a_operand\[5\] MuI.a_operand\[4\] MuI._2866_ vssd1 vssd1
+ vccd1 vccd1 MuI._0809_ sky130_fd_sc_hd__a22o_1
XANTENNA__09199__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _03355_ _03373_ _03372_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a21bo_1
XMuI._4011_ MuI._3109_ MuI._3110_ vssd1 vssd1 vccd1 vccd1 MuI._3111_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _02621_ _05368_ _02619_ _02618_ _02617_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a32o_1
XFILLER_75_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10138__A _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09349__D _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08008__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08008__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6391__A2 MuI._1975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _00279_ _06666_ _00398_ _03378_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08831__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0887__A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5962_ MuI._1787_ MuI._1788_ MuI._1800_ MuI._0769_ vssd1 vssd1 vccd1 vccd1 MuI._1801_
+ sky130_fd_sc_hd__a211o_1
X_11409_ _04094_ _04095_ _04138_ _04139_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nand4_2
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11895__C _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ _05236_ _05237_ _05126_ _05128_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__o211a_1
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4913_ MuI._0440_ MuI._0441_ MuI._0454_ vssd1 vssd1 vccd1 vccd1 MuI._0648_ sky130_fd_sc_hd__a21oi_1
XMuI._5893_ MuI._1721_ MuI._1722_ MuI._1723_ vssd1 vssd1 vccd1 vccd1 MuI._1726_ sky130_fd_sc_hd__and3_1
XFILLER_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13168__B _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4844_ MuI._0560_ MuI._0569_ MuI._0571_ vssd1 vssd1 vccd1 vccd1 MuI._0572_ sky130_fd_sc_hd__o21ai_2
X_06950_ net11 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07166__B _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4775_ MuI._0476_ MuI._0491_ MuI._0494_ vssd1 vssd1 vccd1 vccd1 MuI._0496_ sky130_fd_sc_hd__a21o_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06881_ _04144_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[3\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6514_ MuI._2400_ MuI._2408_ vssd1 vssd1 vccd1 vccd1 MuI._2409_ sky130_fd_sc_hd__and2b_1
XMuI._3726_ MuI.b_operand\[22\] vssd1 vssd1 vccd1 vccd1 MuI._2826_ sky130_fd_sc_hd__buf_2
X_08620_ _01086_ _01085_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__nor2_1
XANTENNA__12400__A2_N _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6445_ MuI._2324_ MuI._2332_ MuI._2322_ vssd1 vssd1 vccd1 vccd1 MuI._2333_ sky130_fd_sc_hd__a21o_1
XMuI._3657_ MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 MuI._2583_ sky130_fd_sc_hd__clkbuf_4
X_08551_ _03400_ _03906_ _01144_ _01149_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__a211oi_1
X_07502_ _00118_ _00119_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__or2_1
XMuI._6376_ MuI._2255_ MuI._2256_ vssd1 vssd1 vccd1 vccd1 MuI._2257_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3588_ MuI._1813_ MuI._0515_ MuI._1329_ vssd1 vssd1 vccd1 vccd1 MuI._1824_ sky130_fd_sc_hd__and3_1
X_08482_ _03099_ _04176_ _04240_ _03056_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4209__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07332__D _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5327_ MuI._1085_ MuI._1086_ MuI._1100_ vssd1 vssd1 vccd1 vccd1 MuI._1103_ sky130_fd_sc_hd__a21o_1
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07433_ _00045_ _00050_ _03002_ _04520_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__and4bb_1
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3968__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3968__B2 MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5258_ MuI._1024_ MuI._1025_ MuI._1026_ vssd1 vssd1 vccd1 vccd1 MuI._1027_ sky130_fd_sc_hd__and3_1
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07364_ _06516_ _05370_ _06489_ _06520_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__a22o_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5765__B MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12043__A2 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4209_ MuI._0768_ MuI._2885_ MuI._3185_ MuI._0559_ vssd1 vssd1 vccd1 vccd1 MuI._3309_
+ sky130_fd_sc_hd__a22oi_1
X_09103_ _06610_ _04122_ _01416_ _01417_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12247__B _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5189_ MuI._0947_ MuI._0948_ MuI._0949_ vssd1 vssd1 vccd1 vccd1 MuI._0951_ sky130_fd_sc_hd__a21o_1
XANTENNA__11251__B1 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07295_ _06588_ _06595_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__and2b_1
XFILLER_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09034_ _03293_ _03895_ _03982_ _03239_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a22oi_2
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07758__B1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1405__B AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ _02325_ _02336_ _02337_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__or3_1
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09867_ _02519_ _02488_ _02489_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__nand3_1
XANTENNA__11857__A2 _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _01431_ _01434_ _01435_ _01415_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07804__B _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13059__A1 _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09798_ _02439_ _02440_ _02436_ _02438_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a211o_1
XANTENNA__13059__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09652__A1_N _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _06622_ _00072_ _00083_ _00414_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__a22oi_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6117__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5659__C MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11760_ _03525_ _04725_ _04432_ _04431_ _04854_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a32o_2
XFILLER_199_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07289__A2 _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _03230_ _03227_ _03229_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a21bo_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _04359_ _04487_ _06428_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__a21oi_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08635__B _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13430_ _01327_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__xor2_4
X_10642_ _03198_ _03201_ _03199_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o21bai_1
XFILLER_41_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3476__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ _06248_ _06249_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__or2b_1
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _03280_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__xnor2_2
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09169__D _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10596__A2 _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12312_ _05042_ _05150_ _05153_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__or3_1
X_13292_ _06199_ _06200_ _06201_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand3_1
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ _03658_ _05047_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__nand2_2
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08370__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1621_ AuI._0693_ AuI._0784_ AuI._0788_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0789_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07267__A _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3923__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _02444_ _02446_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__nand2_1
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11125_ _03874_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__xor2_4
XANTENNA_AuI.pe._726__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1552_ AuI._0661_ AuI._0731_ vssd1 vssd1 vccd1 vccd1 AuI._0732_ sky130_fd_sc_hd__nor2_1
XANTENNA__08961__A2 _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4100__A MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11056_ _02496_ _03801_ _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._1014__A1 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1483_ AuI._0645_ AuI._0651_ AuI._0663_ AuI._0668_ AuI._0634_ vssd1 vssd1 vccd1
+ vccd1 AuI._0669_ sky130_fd_sc_hd__a311o_1
XFILLER_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11848__A2 _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4560_ MuI._0255_ MuI._0202_ MuI._0257_ vssd1 vssd1 vccd1 vccd1 MuI._0259_ sky130_fd_sc_hd__and3_1
X_10007_ _02659_ _02661_ _02660_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a21o_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08098__A _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3511_ MuI._0933_ MuI._0955_ MuI._0966_ vssd1 vssd1 vccd1 vccd1 MuI._0977_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09632__D _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4491_ MuI._0181_ MuI._0182_ vssd1 vssd1 vccd1 vccd1 MuI._0183_ sky130_fd_sc_hd__xor2_1
XFILLER_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__C _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6230_ MuI._2797_ MuI._0438_ vssd1 vssd1 vccd1 vccd1 MuI._2096_ sky130_fd_sc_hd__nand2_1
XMuI._3442_ MuI.a_operand\[27\] MuI.b_operand\[27\] vssd1 vssd1 vccd1 vccd1 MuI._0218_
+ sky130_fd_sc_hd__or2_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11958_ _00216_ _03247_ _05820_ _00217_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__a22o_1
XANTENNA__08826__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6161_ MuI._1483_ MuI._1263_ vssd1 vssd1 vccd1 vccd1 MuI._2020_ sky130_fd_sc_hd__nand2_1
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07730__A _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12993__D _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5939__A2 MuI._0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ _03416_ _03470_ _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a21oi_1
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5112_ MuI._2785_ MuI._2885_ MuI._3185_ MuI._2790_ vssd1 vssd1 vccd1 vccd1 MuI._0866_
+ sky130_fd_sc_hd__a22oi_1
X_11889_ _04662_ _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__and3_1
XFILLER_20_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10794__C _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6092_ MuI._1153_ MuI._2627_ MuI._2914_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._1944_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5043_ MuI._3305_ MuI._0012_ vssd1 vssd1 vccd1 vccd1 MuI._0791_ sky130_fd_sc_hd__or2_1
XFILLER_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4831__A2_N MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ _06056_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__clkbuf_2
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5945_ MuI._0760_ MuI._0761_ MuI._0707_ MuI._0762_ vssd1 vssd1 vccd1 vccd1 MuI._1783_
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__07177__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4127__A1 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._825_ AuI.pe._360_ AuI.pe._362_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[4\]
+ sky130_fd_sc_hd__xor2_1
Xfanout107 net65 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_4
XMuI._5876_ MuI._1631_ MuI._1650_ MuI._1705_ MuI._1706_ vssd1 vssd1 vccd1 vccd1 MuI._1707_
+ sky130_fd_sc_hd__a211o_1
Xfanout118 net46 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_4
XANTENNA__08952__A2 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout129 net25 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_6
X_07982_ _00590_ _00598_ _00599_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__a21boi_2
XANTENNA__12811__A _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._756_ AuI.pe._299_ vssd1 vssd1 vccd1 vccd1 AuI.pe._300_ sky130_fd_sc_hd__inv_2
XFILLER_101_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4827_ MuI.a_operand\[16\] MuI.b_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._0553_
+ sky130_fd_sc_hd__nand2_1
X_09721_ _02348_ _02349_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__and3_1
X_06933_ _04703_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__buf_4
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11839__A2 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._687_ AuI.pe._120_ AuI.pe._004_ AuI.pe._041_ AuI.pe._201_ AuI.pe._234_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._235_ sky130_fd_sc_hd__a221o_1
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4758_ MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 MuI._0477_ sky130_fd_sc_hd__buf_2
XFILLER_110_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11427__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09652_ _06545_ _00303_ _02272_ _02271_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__o2bb2a_1
X_06864_ _03960_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3709_ MuI._2783_ MuI._2784_ MuI._2808_ vssd1 vssd1 vccd1 vccd1 MuI._2809_ sky130_fd_sc_hd__and3_1
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08603_ _06500_ _05025_ _06623_ _06501_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__a22oi_1
XMuI._4689_ MuI._0398_ MuI._0399_ MuI._0400_ vssd1 vssd1 vccd1 vccd1 MuI._0401_ sky130_fd_sc_hd__a21oi_1
X_09583_ _02187_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a21o_1
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06795_ _03217_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__clkbuf_4
XFILLER_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6428_ MuI._2267_ MuI._2312_ MuI._1977_ vssd1 vssd1 vccd1 vccd1 MuI._2314_ sky130_fd_sc_hd__a21oi_1
XANTENNA_AuI.pe._496__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ _00915_ _00930_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._132__138 vssd1 vssd1 vccd1 vccd1 FuI._132__138/HI net138 sky130_fd_sc_hd__conb_1
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08736__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6359_ MuI._2235_ MuI._2236_ MuI._2200_ MuI._2201_ vssd1 vssd1 vccd1 vccd1 MuI._2238_
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _01071_ _01073_ _01072_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07416_ _02948_ _04638_ _00033_ _02894_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__a22oi_1
XFILLER_168_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12016__A2 _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08396_ _01009_ _01013_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07347_ _06643_ _06645_ _06644_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__o21ai_1
XFILLER_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07278_ net38 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12705__B _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ _01540_ _01542_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__or2b_1
XFILLER_164_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07087__A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4986__A1_N MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _02484_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._3877__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11337__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07534__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _03798_ _05391_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__nand2_1
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__C _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _05742_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04614_ _04617_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__nand2_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _02854_ _02868_ _05582_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nand3_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09120__A2 _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _04533_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__xnor2_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11674_ _04466_ _04468_ _04430_ _04222_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o211ai_2
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11215__B1 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ _06325_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._3801__B1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ _03148_ _03147_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__or2b_1
XFILLER_155_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10556_ _03263_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__and2b_1
X_13344_ _06254_ _06255_ _06428_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0983_ AuI._0144_ AuI._0145_ vssd1 vssd1 vccd1 vccd1 AuI._0195_ sky130_fd_sc_hd__and2_1
XFILLER_182_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10487_ _03010_ _03012_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__nand2_1
X_13275_ _06102_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_136_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09187__A2 _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3991_ MuI._2916_ vssd1 vssd1 vccd1 vccd1 MuI._3091_ sky130_fd_sc_hd__clkbuf_4
X_12226_ _05061_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__nand2_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__B _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5730_ MuI._1543_ MuI._1544_ MuI._1052_ MuI._1479_ vssd1 vssd1 vccd1 vccd1 MuI._1546_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12191__A1 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1604_ AuI._0629_ AuI._0644_ AuI._0669_ AuI._0672_ vssd1 vssd1 vccd1 vccd1 AuI._0775_
+ sky130_fd_sc_hd__nand4_1
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12157_ _04853_ _04905_ _04987_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__a211oi_4
XAuI.pe._610_ AuI.pe._055_ AuI.pe._133_ AuI.pe._150_ AuI.pe._029_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._163_ sky130_fd_sc_hd__a22o_1
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__A _02801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5661_ MuI._1468_ MuI._1469_ vssd1 vssd1 vccd1 vccd1 MuI._1470_ sky130_fd_sc_hd__nand2_1
X_11108_ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__inv_2
XAuI._1535_ AuI._0717_ AuI._0658_ vssd1 vssd1 vccd1 vccd1 AuI._0718_ sky130_fd_sc_hd__xor2_1
X_12088_ _04773_ _04775_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__nand2_1
XAuI.pe._541_ AuI.pe._062_ AuI.pe._050_ AuI.pe._042_ AuI.pe._072_ AuI.pe._098_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._099_ sky130_fd_sc_hd__a221o_1
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4612_ MuI._2826_ MuI.b_operand\[21\] MuI._0315_ vssd1 vssd1 vccd1 vccd1 MuI._0316_
+ sky130_fd_sc_hd__and3_1
XMuI._5592_ MuI._1377_ MuI._1378_ MuI._1392_ vssd1 vssd1 vccd1 vccd1 MuI._1394_ sky130_fd_sc_hd__a21oi_1
X_11039_ _03783_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1466_ AuI._0346_ AuI._0342_ vssd1 vssd1 vccd1 vccd1 AuI._0652_ sky130_fd_sc_hd__or2b_1
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._472_ AuI.pe._035_ vssd1 vssd1 vccd1 vccd1 AuI.pe._036_ sky130_fd_sc_hd__buf_2
XMuI._4543_ MuI._0239_ vssd1 vssd1 vccd1 vccd1 MuI._0241_ sky130_fd_sc_hd__inv_2
XFILLER_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1397_ AuI._0258_ AuI._0584_ AuI._0585_ AuI._0586_ vssd1 vssd1 vccd1 vccd1 AuI._0587_
+ sky130_fd_sc_hd__and4_1
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4474_ MuI._0024_ MuI._0026_ vssd1 vssd1 vccd1 vccd1 MuI._0165_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6213_ MuI._2035_ MuI._2037_ MuI._2036_ vssd1 vssd1 vccd1 vccd1 MuI._2078_ sky130_fd_sc_hd__o21ai_1
XFILLER_206_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3425_ MuI.a_operand\[28\] MuI.a_operand\[27\] MuI.a_operand\[29\] MuI.a_operand\[30\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0032_ sky130_fd_sc_hd__and4_1
XFILLER_45_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11454__B1 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1171__A0 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6144_ MuI._2001_ vssd1 vssd1 vccd1 vccd1 MuI._2002_ sky130_fd_sc_hd__inv_2
X_08250_ _00857_ _00862_ _00866_ _00867_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__o211ai_4
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__A2 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08870__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07201_ _06500_ _06476_ _06489_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__a22oi_1
XMuI._6075_ MuI._1885_ MuI._1900_ MuI._1925_ vssd1 vssd1 vccd1 vccd1 MuI._1926_ sky130_fd_sc_hd__o21ai_1
XFILLER_193_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5793__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08181_ _00393_ _00405_ _00392_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._4005__A MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11132__D _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5026_ MuI._0653_ MuI._0770_ MuI._0769_ MuI._0765_ vssd1 vssd1 vccd1 vccd1 MuI._0772_
+ sky130_fd_sc_hd__a211o_1
XFILLER_146_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__A1 _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07132_ _04100_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11710__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6337__A2 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__A _00610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06804__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07063_ _06098_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_173_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5928_ MuI._1556_ MuI._1643_ MuI._1641_ vssd1 vssd1 vccd1 vccd1 MuI._1764_ sky130_fd_sc_hd__a21o_1
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12541__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._808_ AuI.pe.significand\[13\] AuI.pe.significand\[14\] AuI.pe.significand\[15\]
+ AuI.pe._367_ vssd1 vssd1 vccd1 vccd1 AuI.pe._347_ sky130_fd_sc_hd__or4_1
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5859_ MuI._0750_ MuI._1686_ MuI._1685_ vssd1 vssd1 vccd1 vccd1 MuI._1688_ sky130_fd_sc_hd__a21o_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07965_ _00277_ _00582_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__or2_1
XANTENNA__08138__B1 _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._739_ AuI.pe._106_ AuI.pe._150_ AuI.pe._280_ AuI.pe._282_ AuI.pe._283_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._284_ sky130_fd_sc_hd__a2111o_1
X_09704_ _02301_ _02293_ _02300_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__nand3_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06916_ _04520_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__buf_6
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4394__B MuI._0076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07896_ _00505_ _00513_ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09635_ _02271_ _02273_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__nor2_1
XFILLER_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06847_ _03777_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[30\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07361__A1 _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06778_ _03035_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[17\] sky130_fd_sc_hd__clkbuf_1
X_09566_ _06494_ _06495_ _00082_ _00084_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__and4_1
XFILLER_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08466__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _01066_ _01119_ _01133_ _01134_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__a211oi_2
XFILLER_169_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09497_ _01978_ _01970_ _01977_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__nand3_1
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10799__A2 _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07664__A2 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ _01017_ _01050_ _01064_ _01065_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__o211ai_4
XANTENNA__10089__A_N _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08379_ _00978_ _00979_ _00980_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__o21bai_1
XFILLER_184_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._083_ FuI._047_ vssd1 vssd1 vccd1 vccd1 FuI._016_ sky130_fd_sc_hd__clkbuf_1
X_10410_ _03004_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__xnor2_2
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11390_ _02757_ _04017_ _01988_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__o21a_1
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07416__A2 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06714__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _03030_ _03031_ _03032_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a21o_1
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10236__A _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _02815_ _05883_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__o21a_1
X_10272_ _00683_ _00682_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__or2b_1
XFILLER_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07248__C _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12011_ _04683_ _04691_ _04690_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21o_1
XANTENNA__08377__B1 _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07545__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1320_ AuI._0486_ AuI._0490_ AuI._0501_ AuI._0516_ vssd1 vssd1 vccd1 vccd1 AuI._0517_
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12913_ _05695_ _05707_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__and2b_1
XAuI._1251_ AuI._0448_ AuI._0451_ vssd1 vssd1 vccd1 vccd1 AuI._0453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6264__A1 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07352__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07352__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12844_ _05714_ _05715_ _05725_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__and3_1
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1182_ AuI._0263_ AuI._0383_ AuI._0387_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0388_
+ sky130_fd_sc_hd__a211o_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08376__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07280__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05610_ _05651_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or3_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1153__A0 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4190_ MuI._3287_ MuI._3289_ vssd1 vssd1 vccd1 vccd1 MuI._3290_ sky130_fd_sc_hd__xor2_1
XFILLER_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _04522_ _04523_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__nand3_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__D _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11657_ _02983_ _02984_ _04972_ _00421_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__nand4_1
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _03993_ _02216_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2b_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11588_ _04374_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nor2_1
XFILLER_183_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08542__C _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _06226_ _06176_ _06236_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__and3_1
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10539_ net25 vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__clkbuf_4
XAuI._0966_ AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0178_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._6040__A MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09357__D net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6831_ MuI._2698_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2747_ sky130_fd_sc_hd__and2b_1
XANTENNA__08261__D _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13258_ _06112_ _06114_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__nand2_1
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0895__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07158__C net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0897_ AuI._0115_ AuI._0116_ vssd1 vssd1 vccd1 vccd1 AuI._0117_ sky130_fd_sc_hd__or2_2
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6762_ MuI._2588_ MuI._2597_ MuI._2601_ vssd1 vssd1 vccd1 vccd1 MuI._2681_ sky130_fd_sc_hd__and3_1
XMuI._3974_ MuI._2971_ MuI._2969_ MuI._2970_ vssd1 vssd1 vccd1 vccd1 MuI._3074_ sky130_fd_sc_hd__a21o_1
X_12209_ _03024_ _05831_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nand2_1
XFILLER_151_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13189_ _02841_ _06011_ _02839_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__a21o_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5713_ MuI._2852_ MuI.a_operand\[15\] MuI._0017_ MuI._3396_ vssd1 vssd1 vccd1
+ vccd1 MuI._1528_ sky130_fd_sc_hd__and4_1
XFILLER_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0967__A0 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6693_ MuI._2002_ MuI._2602_ vssd1 vssd1 vccd1 vccd1 MuI._2606_ sky130_fd_sc_hd__or2_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1503__B AuI._0586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5644_ MuI._1408_ MuI._1447_ MuI._1449_ MuI._1451_ vssd1 vssd1 vccd1 vccd1 MuI._1452_
+ sky130_fd_sc_hd__a31o_1
XAuI._1518_ AuI._0702_ vssd1 vssd1 vccd1 vccd1 AuI._0703_ sky130_fd_sc_hd__buf_2
XFILLER_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07750_ _00334_ _00339_ _00366_ _00367_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._3830__C MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._524_ AuI.pe._075_ AuI.pe._083_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[6\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_84_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5575_ MuI._1341_ MuI._1375_ vssd1 vssd1 vccd1 vccd1 MuI._1376_ sky130_fd_sc_hd__xor2_2
X_06701_ _02205_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07681_ net50 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__buf_2
XAuI._1449_ AuI._0422_ AuI._0439_ AuI._0444_ vssd1 vssd1 vccd1 vccd1 AuI._0635_ sky130_fd_sc_hd__and3_1
XFILLER_53_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._455_ AuI.pe._005_ AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 AuI.pe._021_ sky130_fd_sc_hd__and2b_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4526_ MuI._0213_ MuI._0221_ vssd1 vssd1 vccd1 vccd1 MuI._0222_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09420_ _01962_ _02039_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__and2b_1
XFILLER_52_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07902__B _00519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07190__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4457_ MuI._0139_ MuI._0144_ MuI._0015_ vssd1 vssd1 vccd1 vccd1 MuI._0146_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08717__C _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _06544_ _04445_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__nand2_1
XFILLER_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07621__C _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5757__C MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _00262_ _00272_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__nand2_1
XMuI._4388_ MuI._0059_ MuI._0063_ MuI._0069_ MuI._0070_ vssd1 vssd1 vccd1 vccd1 MuI._0071_
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _06583_ _00287_ _00267_ _02593_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22oi_2
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6127_ MuI._3147_ MuI._1902_ MuI._1982_ vssd1 vssd1 vccd1 vccd1 MuI._1983_ sky130_fd_sc_hd__o21a_1
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08233_ _00548_ _00850_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._5766__B1 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout130_A net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6058_ MuI._1904_ MuI._1906_ vssd1 vssd1 vccd1 vccd1 MuI._1907_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _02377_ _05702_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__nand2_1
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5009_ MuI._0751_ MuI._0752_ vssd1 vssd1 vccd1 vccd1 MuI._0753_ sky130_fd_sc_hd__nand2_1
X_07115_ _06421_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[26\] sky130_fd_sc_hd__clkbuf_2
XFILLER_109_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _00455_ _00472_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__nor2_2
XANTENNA__10056__A _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07046_ _05917_ _02042_ _02151_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__and3_1
XFILLER_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13352__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__B _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12271__A _05092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0958__A0 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07365__A _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09283__C _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5297__A2 MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08997_ _01612_ _01611_ _01613_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__nor4b_1
XANTENNA__07582__A1 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07948_ _00012_ _00040_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__and2_4
XANTENNA_AuI.pe._603__A1_N AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._138__144 vssd1 vssd1 vccd1 vccd1 FuI._138__144/HI net144 sky130_fd_sc_hd__conb_1
XANTENNA__12458__A2 _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5049__A2 MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6246__A1 MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _00350_ _00353_ _00495_ _00496_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a211oi_1
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09618_ _02238_ _02239_ _02252_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10890_ _02485_ _00785_ _03082_ _06565_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a22o_1
XFILLER_55_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06709__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__inv_2
XANTENNA__09087__A1 _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11969__A1 _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__B2 _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3468__B MuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _05196_ _05199_ _05322_ _05323_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__o211a_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11511_ _04253_ _04254_ _04291_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__o211ai_4
XFILLER_200_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12446__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12491_ _05346_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__nor2_1
XFILLER_184_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._135_ FuI._019_ net141 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[6\] sky130_fd_sc_hd__dlxtn_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11350__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ _04217_ _04200_ _04201_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__and3_1
XFILLER_184_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._066_ FuI.a_operand\[28\] FuI.a_operand\[29\] net105 vssd1 vssd1 vccd1 vccd1
+ FuI._034_ sky130_fd_sc_hd__o21a_1
XANTENNA__08598__B1 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__C net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0820_ AuI._0038_ net15 AuI._0039_ net14 vssd1 vssd1 vccd1 vccd1 AuI._0040_ sky130_fd_sc_hd__a22o_1
XFILLER_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ _04142_ _04143_ _03902_ _03904_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__o211a_1
XFILLER_180_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13112_ _02841_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nand2_1
X_10324_ _03007_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__nand3_1
XANTENNA_input60_A b_operand[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._409__B_N AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4732__A1 MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10255_ _02727_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09474__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13043_ _05911_ _05913_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nand2_1
XFILLER_106_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10186_ _03110_ _05209_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__and2b_1
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3690_ MuI.a_operand\[10\] vssd1 vssd1 vccd1 vccd1 MuI._2790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6019__B MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1303_ AuI._0498_ AuI._0499_ AuI._0500_ vssd1 vssd1 vccd1 vccd1 AuI._0501_ sky130_fd_sc_hd__or3_2
XFILLER_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1374__A0 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5360_ MuI._1122_ MuI._1123_ MuI._1138_ vssd1 vssd1 vccd1 vccd1 MuI._1139_ sky130_fd_sc_hd__nand3_1
XFILLER_74_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1234_ AuI._0256_ vssd1 vssd1 vccd1 vccd1 AuI._0437_ sky130_fd_sc_hd__buf_2
XFILLER_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4311_ MuI._3408_ MuI._3410_ vssd1 vssd1 vccd1 vccd1 MuI._3411_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5291_ MuI._2975_ MuI._2976_ MuI._0245_ MuI._0321_ vssd1 vssd1 vccd1 vccd1 MuI._1063_
+ sky130_fd_sc_hd__and4_1
X_12827_ _05695_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1165_ AuI._0263_ AuI._0371_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0372_ sky130_fd_sc_hd__a21oi_2
XFILLER_188_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4242_ MuI._2796_ MuI._2791_ vssd1 vssd1 vccd1 vccd1 MuI._3342_ sky130_fd_sc_hd__nand2_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__B1 _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08825__A1 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ _06439_ _05391_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nand2_1
XAuI._1096_ AuI._0209_ AuI._0305_ vssd1 vssd1 vccd1 vccd1 AuI._0306_ sky130_fd_sc_hd__or2_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08825__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5296__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4173_ MuI._3270_ MuI._3272_ vssd1 vssd1 vccd1 vccd1 MuI._3273_ sky130_fd_sc_hd__or2_1
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11709_ _02669_ _05906_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__nand2_1
XFILLER_187_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _05557_ _05558_ _05471_ _05473_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a211o_1
XFILLER_175_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08589__B1 _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4971__A1 MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4971__B2 MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07169__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._577__A AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0949_ AuI._0110_ AuI._0160_ vssd1 vssd1 vccd1 vccd1 AuI._0161_ sky130_fd_sc_hd__and2b_1
XFILLER_171_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6814_ MuI.Exception MuI._2731_ MuI._2733_ vssd1 vssd1 vccd1 vccd1 MuI._2737_
+ sky130_fd_sc_hd__nor3_2
X_08920_ _01534_ _01536_ _01535_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a21o_1
XFILLER_131_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3957_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._2876_ vssd1 vssd1 vccd1
+ vccd1 MuI._3057_ sky130_fd_sc_hd__o31a_1
XMuI._6745_ MuI._2476_ MuI._1747_ vssd1 vssd1 vccd1 vccd1 MuI._2663_ sky130_fd_sc_hd__nor2_1
XANTENNA__07185__A _06470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _01447_ _01448_ _01453_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a21o_1
XANTENNA__11896__B1 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6676_ MuI._2579_ MuI._2586_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2587_ sky130_fd_sc_hd__mux2_1
X_07802_ _00416_ _00417_ _00418_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a21o_1
XANTENNA__12241__D _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3888_ MuI._2981_ MuI._2982_ MuI._2987_ vssd1 vssd1 vccd1 vccd1 MuI._2988_ sky130_fd_sc_hd__nand3_1
XFILLER_85_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08782_ _01396_ _01399_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5627_ MuI._1376_ MuI._1432_ vssd1 vssd1 vccd1 vccd1 MuI._1433_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07733_ _03497_ _04122_ _00323_ _00322_ vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__a31o_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._507_ AuI.pe._033_ AuI.pe._050_ AuI.pe._042_ AuI.pe._045_ AuI.pe._067_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._068_ sky130_fd_sc_hd__a221o_1
XFILLER_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5558_ MuI._1347_ MuI._1355_ MuI._1356_ vssd1 vssd1 vccd1 vccd1 MuI._1357_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07664_ _03443_ _06446_ _04111_ _00281_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a22oi_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12860__A2 _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4509_ MuI._0200_ MuI._0201_ MuI._0191_ MuI._0195_ vssd1 vssd1 vccd1 vccd1 MuI._0203_
+ sky130_fd_sc_hd__o211ai_1
XAuI.pe._438_ AuI.pe.significand\[23\] AuI.pe.significand\[24\] vssd1 vssd1 vccd1
+ vccd1 AuI.pe._005_ sky130_fd_sc_hd__and2b_1
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _01919_ _01920_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__or2_1
XFILLER_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5489_ MuI._1217_ MuI._1226_ MuI._1225_ vssd1 vssd1 vccd1 vccd1 MuI._1281_ sky130_fd_sc_hd__a21o_1
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11154__B _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _00211_ _00210_ _00025_ _06676_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__a211o_1
XANTENNA__07351__C _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09334_ _01946_ _01950_ _01951_ _01835_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__o211ai_2
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12612__A2 _05476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10623__A1 _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _01842_ _01841_ _01810_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a21o_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__A2 _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ _00632_ _00629_ _00631_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__a21o_1
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ _01813_ _01770_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _00762_ _00763_ _00755_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__a21o_1
XFILLER_20_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08078_ _00292_ _00259_ _00694_ _00695_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a22o_1
XFILLER_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07029_ _05735_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[27\] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07807__B _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07095__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ _06023_ _02709_ _02064_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__or3b_1
XFILLER_103_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10233__B _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._532__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ _04768_ _04769_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand4_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1356__A0 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07542__B _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10942_ _03489_ _03672_ _03673_ _03679_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__a31o_1
XFILLER_84_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08357__C _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ _02658_ _05638_ _00163_ _02593_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__a22oi_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _05475_ _05476_ _05301_ _05306_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__o211a_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08807__A1 _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08807__B2 _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5694__A MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ _00270_ _05649_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__nand2_1
XFILLER_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._599__A1 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._599__B2 AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ _05326_ _05328_ _05178_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__o21ai_2
XFuI._118_ FuI._050_ FuI._056_ FuI._024_ FuI._029_ FuI.a_operand\[15\] vssd1 vssd1
+ vccd1 vccd1 FuI._005_ sky130_fd_sc_hd__o311a_1
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12367__A1 _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11425_ _04196_ _04198_ _04199_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__a21o_1
XFILLER_153_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12904__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _04115_ _04125_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and3_1
XANTENNA__06902__A _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4860_ MuI._0572_ MuI._0585_ MuI._0586_ MuI._0587_ vssd1 vssd1 vccd1 vccd1 MuI._0589_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12119__B2 _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__C net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _02994_ _02995_ _00698_ _00702_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__o211a_1
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11287_ _03943_ _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__and3_1
XMuI._3811_ MuI._2907_ MuI._2910_ vssd1 vssd1 vccd1 vccd1 MuI._2911_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12342__C _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4791_ MuI._0462_ MuI._0512_ vssd1 vssd1 vccd1 vccd1 MuI._0513_ sky130_fd_sc_hd__nor2_1
X_13026_ _05752_ _05920_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10238_ _02918_ _02922_ _02814_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__o21bai_1
XANTENNA__11239__B _04000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6530_ MuI._2419_ MuI._2425_ vssd1 vssd1 vccd1 vccd1 MuI._2426_ sky130_fd_sc_hd__and2_1
XANTENNA__10143__B _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3742_ MuI._2840_ MuI._2841_ vssd1 vssd1 vccd1 vccd1 MuI._2842_ sky130_fd_sc_hd__nand2_1
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _02845_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nand2_2
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07155__D _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6461_ MuI._2320_ MuI._2327_ vssd1 vssd1 vccd1 vccd1 MuI._2350_ sky130_fd_sc_hd__nand2_1
XFILLER_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3673_ MuI._2572_ MuI._2736_ MuI._2743_ vssd1 vssd1 vccd1 vccd1 MuI._2748_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI.pe._523__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5412_ MuI.a_operand\[7\] MuI.a_operand\[6\] MuI._3402_ MuI._3396_ vssd1 vssd1
+ vccd1 vccd1 MuI._1196_ sky130_fd_sc_hd__and4_1
XANTENNA__12062__A2_N _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1347__A0 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6392_ MuI._2269_ MuI._2270_ MuI._2100_ MuI._2273_ vssd1 vssd1 vccd1 vccd1 MuI._2274_
+ sky130_fd_sc_hd__and4b_1
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10302__B1 _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4492__B MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3692__B2 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5343_ MuI._1110_ MuI._1112_ vssd1 vssd1 vccd1 vccd1 MuI._1121_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1217_ AuI._0288_ AuI._0249_ vssd1 vssd1 vccd1 vccd1 AuI._0421_ sky130_fd_sc_hd__nor2_1
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5274_ MuI._1041_ MuI._1042_ MuI._1037_ vssd1 vssd1 vccd1 vccd1 MuI._1045_ sky130_fd_sc_hd__a21o_1
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07380_ _06680_ _05112_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__and2_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1148_ AuI._0274_ AuI._0188_ AuI._0355_ vssd1 vssd1 vccd1 vccd1 AuI._0356_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4225_ MuI._3315_ MuI._3322_ MuI._3324_ vssd1 vssd1 vccd1 vccd1 MuI._3325_ sky130_fd_sc_hd__a21o_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1509__A AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1079_ AuI._0171_ AuI._0182_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0290_ sky130_fd_sc_hd__mux2_1
XMuI._4156_ MuI._3211_ MuI._3197_ vssd1 vssd1 vccd1 vccd1 MuI._3256_ sky130_fd_sc_hd__nand2_1
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09050_ _01208_ _01579_ _01581_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__o31a_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ _00339_ _00587_ _00586_ _00564_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a211oi_1
XMuI._4087_ MuI._0801_ MuI._2967_ MuI._3184_ MuI._3186_ vssd1 vssd1 vccd1 vccd1 MuI._3187_
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06812__A _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__B _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ _02341_ _02340_ _02603_ _02610_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XFILLER_132_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _01518_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__xor2_1
XMuI._4989_ MuI._0727_ MuI._0729_ vssd1 vssd1 vccd1 vccd1 MuI._0731_ sky130_fd_sc_hd__nor2_1
XANTENNA__11869__B1 _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _02538_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nor2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6728_ MuI._2464_ MuI._2637_ vssd1 vssd1 vccd1 vccd1 MuI._2644_ sky130_fd_sc_hd__or2_1
XFILLER_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08834_ _01450_ _01451_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__nor2_1
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6659_ MuI._2505_ MuI._2509_ MuI._2559_ MuI._2563_ MuI._2567_ vssd1 vssd1 vccd1
+ vccd1 MuI._2568_ sky130_fd_sc_hd__o2111a_1
XFILLER_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08765_ _03002_ _06443_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__nand2_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _00298_ _00317_ _00332_ _00333_ vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__a211o_1
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13491__C1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ _01311_ _01312_ _01313_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__nor3_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ _00261_ _00264_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__and2b_1
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ _00192_ _00193_ _00194_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__a21o_1
XFILLER_201_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _01929_ _01930_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a21o_1
XFILLER_167_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06706__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _01644_ _01851_ _01864_ _01865_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__o211a_1
XFILLER_167_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__xor2_1
XFILLER_182_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6137__B1 MuI._1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _03152_ _06623_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__and2_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11021__A1 _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _02862_ _04865_ _02745_ _02719_ _04929_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a32o_1
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06722__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _03891_ _03892_ _03881_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09455__D _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10780__B1 _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 ALU_Output[17] sky130_fd_sc_hd__buf_2
X_11072_ _03645_ _03643_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__and2b_1
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 ALU_Output[27] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 ALU_Output[8] sky130_fd_sc_hd__buf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10023_ _02687_ _02688_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__nor3_1
XANTENNA__08725__B1 _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input23_A a_operand[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5112__B2 MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _04790_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nand2_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._680__A AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _03331_ _03484_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_1
XFILLER_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0937__B_N AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1002_ net41 net9 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0214_ sky130_fd_sc_hd__mux2_1
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10856_ _03585_ _03586_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__or2b_1
XFILLER_204_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09199__B _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4010_ MuI._3014_ MuI._3016_ MuI._3013_ vssd1 vssd1 vccd1 vccd1 MuI._3110_ sky130_fd_sc_hd__o21ba_1
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _03337_ _03376_ _03512_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__o21ai_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12526_ _05381_ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__or2_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10138__B _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12457_ _00077_ _05520_ _05161_ _05160_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__a31o_1
XANTENNA__08008__A2 _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08831__B _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output91_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5961_ MuI._0737_ MuI._0767_ MuI._1799_ vssd1 vssd1 vccd1 vccd1 MuI._1800_ sky130_fd_sc_hd__a21oi_1
X_11408_ _04107_ _04109_ _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__o21ba_1
XFILLER_172_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12388_ _05232_ _05233_ _05235_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4912_ MuI._0632_ MuI._0634_ MuI._0645_ vssd1 vssd1 vccd1 vccd1 MuI._0646_ sky130_fd_sc_hd__and3_1
XMuI._5892_ MuI._1721_ MuI._1722_ MuI._1723_ vssd1 vssd1 vccd1 vccd1 MuI._1724_ sky130_fd_sc_hd__a21oi_2
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11339_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__and2_1
XANTENNA__10154__A _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4843_ MuI._0511_ MuI._0513_ vssd1 vssd1 vccd1 vccd1 MuI._0571_ sky130_fd_sc_hd__xor2_1
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08716__B1 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3901__A2 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4774_ MuI._0476_ MuI._0491_ MuI._0494_ vssd1 vssd1 vccd1 vccd1 MuI._0495_ sky130_fd_sc_hd__nand3_1
XANTENNA__13465__A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _05900_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06880_ _04133_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__and3_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3725_ MuI._0614_ MuI._2385_ MuI._2330_ MuI._0361_ vssd1 vssd1 vccd1 vccd1 MuI._2825_
+ sky130_fd_sc_hd__a22oi_1
XMuI._6513_ MuI._2405_ MuI._2406_ vssd1 vssd1 vccd1 vccd1 MuI._2408_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07463__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1511__B AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09381__C net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3656_ MuI._2462_ MuI._2506_ MuI._2561_ vssd1 vssd1 vccd1 vccd1 MuI._2572_ sky130_fd_sc_hd__or3_1
XMuI._6444_ MuI._2325_ vssd1 vssd1 vccd1 vccd1 MuI._2332_ sky130_fd_sc_hd__inv_2
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08550_ _01166_ _01167_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__and2_1
XFILLER_208_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6375_ MuI._1942_ MuI._1944_ MuI._1943_ vssd1 vssd1 vccd1 vccd1 MuI._2256_ sky130_fd_sc_hd__o21ba_1
X_07501_ _00115_ _00117_ _00116_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__a21oi_1
XMuI._3587_ MuI._1802_ vssd1 vssd1 vccd1 vccd1 MuI._1813_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08481_ _00095_ _00096_ _00271_ _04229_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._4008__A MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5326_ MuI._1074_ MuI._1078_ vssd1 vssd1 vccd1 vccd1 MuI._1102_ sky130_fd_sc_hd__xor2_1
XANTENNA__12809__A _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07432_ _00046_ _00047_ _00048_ _00049_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a22oi_2
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06807__A _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5257_ MuI._2871_ MuI._2330_ MuI._0901_ MuI._0898_ vssd1 vssd1 vccd1 vccd1 MuI._1026_
+ sky130_fd_sc_hd__a31o_1
XFILLER_149_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3968__A2 MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3847__A MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ _06663_ _05316_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5765__C MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4208_ MuI._0559_ MuI.a_operand\[20\] MuI._3306_ MuI._3307_ vssd1 vssd1 vccd1
+ vccd1 MuI._3308_ sky130_fd_sc_hd__and4_1
XANTENNA__13240__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ _01713_ _01718_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__xor2_1
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5188_ MuI._0947_ MuI._0948_ MuI._0949_ vssd1 vssd1 vccd1 vccd1 MuI._0950_ sky130_fd_sc_hd__nand3_1
XANTENNA__11251__A1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07294_ _06592_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nor2_1
XFILLER_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4139_ MuI._3237_ MuI._3238_ MuI._2817_ MuI._2330_ vssd1 vssd1 vccd1 vccd1 MuI._3239_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09033_ _01649_ _01647_ _01648_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nand3_1
XANTENNA__08741__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11003__A1 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10064__A _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _02037_ _02594_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__or2b_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _02488_ _02489_ _02519_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a21o_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09380__B1 _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08817_ _01413_ _01414_ _01365_ _01381_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__o211a_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _02406_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__inv_2
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13059__A2 _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _02582_ _02647_ _00089_ _00082_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__and4_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6117__B MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5659__D MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _00986_ _00987_ _01002_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__and3_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10710_ _03428_ _03426_ _03427_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__nand3_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _04485_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nor2_1
XFILLER_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06717__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08635__C _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _03202_ _03210_ _03209_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a21o_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11342__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A2 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07446__B1 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ _06225_ _06247_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or2b_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10572_ _03004_ _03107_ _03281_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a21oi_2
XFILLER_194_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12311_ _05042_ _05150_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ _06061_ _06137_ _06138_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o21ai_2
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _05078_ _05079_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nor2_2
XFILLER_182_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3592__B1 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3492__A MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08370__C net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1620_ AuI._0617_ AuI._0787_ vssd1 vssd1 vccd1 vccd1 AuI._0788_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ _02581_ _04881_ _02447_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__o21ai_1
XFILLER_123_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1551_ AuI._0727_ AuI._0650_ vssd1 vssd1 vccd1 vccd1 AuI._0731_ sky130_fd_sc_hd__and2b_1
X_11124_ _03705_ _03707_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__a21oi_4
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4100__B MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1482_ AuI._0664_ AuI._0666_ AuI._0667_ vssd1 vssd1 vccd1 vccd1 AuI._0668_ sky130_fd_sc_hd__or3b_1
X_11055_ _02485_ _03082_ _00789_ _06565_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a22o_1
XFILLER_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09371__B1 _01891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _02672_ _02671_ _02673_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__nor3_2
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5097__B1 MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3510_ MuI._0911_ MuI._0922_ vssd1 vssd1 vccd1 vccd1 MuI._0966_ sky130_fd_sc_hd__nor2_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__B _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4490_ MuI._0037_ MuI._0047_ vssd1 vssd1 vccd1 vccd1 MuI._0182_ sky130_fd_sc_hd__xnor2_2
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07433__D _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3441_ MuI._0163_ MuI._0185_ MuI._0196_ vssd1 vssd1 vccd1 vccd1 MuI._0207_ sky130_fd_sc_hd__a21bo_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _02905_ _02959_ _05767_ _05820_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nand4_1
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6160_ MuI._0779_ MuI._1010_ MuI._3000_ MuI._2754_ vssd1 vssd1 vccd1 vccd1 MuI._2019_
+ sky130_fd_sc_hd__and4_1
XANTENNA__08826__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _03469_ _03467_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__and2b_1
XANTENNA__07730__B _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5111_ MuI._0858_ MuI._0863_ MuI._0864_ vssd1 vssd1 vccd1 vccd1 MuI._0865_ sky130_fd_sc_hd__a21bo_1
X_11888_ _04696_ _04697_ _04525_ _04546_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o211ai_1
XFILLER_177_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6091_ MuI._0735_ MuI._2813_ MuI._2627_ MuI._2682_ vssd1 vssd1 vccd1 vccd1 MuI._1943_
+ sky130_fd_sc_hd__and4_1
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10794__D _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ _03567_ _03565_ _03566_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand3_1
XFILLER_186_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10149__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5042_ MuI._0146_ MuI._0787_ MuI._3304_ MuI._0013_ MuI._0788_ vssd1 vssd1 vccd1
+ vccd1 MuI._0789_ sky130_fd_sc_hd__o2111a_1
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0898__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07988__A1 _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ _02970_ _02724_ _05362_ _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a211o_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ _06355_ _06357_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__and2b_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12083__B _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5944_ MuI._1779_ MuI._1781_ vssd1 vssd1 vccd1 vccd1 MuI._1782_ sky130_fd_sc_hd__or2_1
XFILLER_114_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07177__B _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._824_ AuI.pe._330_ AuI.pe._341_ AuI.pe._358_ AuI.pe._361_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._362_ sky130_fd_sc_hd__a31o_1
XANTENNA__11941__C1 _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net64 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_6
XMuI._5875_ MuI._1702_ MuI._1704_ MuI._1667_ vssd1 vssd1 vccd1 vccd1 MuI._1706_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout119 net45 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_6
X_07981_ _00260_ _00597_ _00591_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__or3_1
XFILLER_141_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._755_ AuI.pe._373_ AuI.pe._379_ AuI.pe._298_ vssd1 vssd1 vccd1 vccd1 AuI.pe._299_
+ sky130_fd_sc_hd__or3_1
XANTENNA__12811__B _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4826_ MuI.a_operand\[18\] MuI.a_operand\[17\] MuI.b_operand\[1\] MuI.b_operand\[0\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0552_ sky130_fd_sc_hd__and4_1
X_09720_ _02355_ _02363_ _02364_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a21bo_1
XFILLER_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06932_ net8 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4945__B MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._686_ AuI.pe._385_ AuI.pe._025_ AuI.pe._022_ AuI.pe._211_ AuI.pe._036_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._234_ sky130_fd_sc_hd__a221o_1
XANTENNA__07193__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4757_ MuI._0465_ MuI._0473_ MuI._0475_ vssd1 vssd1 vccd1 vccd1 MuI._0476_ sky130_fd_sc_hd__a21o_1
X_09651_ _02251_ _02250_ _02242_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21o_1
XANTENNA__11427__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06863_ net132 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3708_ MuI._2794_ MuI._2806_ MuI._2807_ vssd1 vssd1 vccd1 vccd1 MuI._2808_ sky130_fd_sc_hd__a21bo_1
X_08602_ net108 _04961_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__nand2_1
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4688_ MuI._0397_ MuI._0396_ vssd1 vssd1 vccd1 vccd1 MuI._0400_ sky130_fd_sc_hd__and2b_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _02211_ _02214_ _02143_ _02188_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__o211a_1
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06794_ net50 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__buf_2
XMuI._6427_ MuI._1977_ MuI._2267_ MuI._2312_ vssd1 vssd1 vccd1 vccd1 MuI._2313_ sky130_fd_sc_hd__and3_1
XMuI._3639_ MuI._2374_ vssd1 vssd1 vccd1 vccd1 MuI._2385_ sky130_fd_sc_hd__buf_2
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ _01143_ _01150_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__nand2_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08736__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6358_ MuI._2200_ MuI._2201_ MuI._2235_ MuI._2236_ vssd1 vssd1 vccd1 vccd1 MuI._2237_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_51_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08464_ _00221_ _04251_ _01081_ _01079_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a31o_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5309_ MuI._1081_ MuI._1082_ vssd1 vssd1 vccd1 vccd1 MuI._1083_ sky130_fd_sc_hd__nor2_1
XMuI._6289_ MuI._2138_ MuI._2137_ vssd1 vssd1 vccd1 vccd1 MuI._2161_ sky130_fd_sc_hd__and2b_1
X_07415_ _00032_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__buf_4
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _01010_ _01012_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07346_ _06536_ _06538_ _06535_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__o21bai_1
XFILLER_176_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3727__D MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5792__A MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ net68 vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__clkbuf_4
XFILLER_191_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ _01556_ _01558_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__and2_1
XFILLER_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07600__B1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _02576_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__or2_1
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3877__A1 MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3877__B2 MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__A _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12440__C _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__inv_2
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11337__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5079__B1 MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__D _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ _03842_ _05273_ _05643_ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a31oi_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07831__A _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ _04322_ _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o21a_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _05667_ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21a_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__nor2_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _04430_ _04222_ _04466_ _04468_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a211o_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11215__A1 _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ _03842_ _05853_ _06281_ _06279_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a31o_1
X_10624_ _03181_ _03218_ _03215_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o21ai_2
XANTENNA_MuI._3801__A1 MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__B2 _03974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3801__B2 MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__A1 _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13343_ _06196_ _06204_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__nand2_1
X_10555_ _00791_ _03090_ _03262_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__or3_1
XAuI._0982_ AuI._0141_ AuI._0142_ vssd1 vssd1 vccd1 vccd1 AuI._0194_ sky130_fd_sc_hd__and2_1
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07278__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ _06182_ _06183_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _03187_ _03188_ _03182_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a21o_1
XFILLER_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3990_ MuI._2999_ MuI._3002_ vssd1 vssd1 vccd1 vccd1 MuI._3090_ sky130_fd_sc_hd__nand2_1
XFILLER_182_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _05060_ _05059_ _05057_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._4463__A1_N MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1603_ AuI._0259_ AuI._0773_ AuI._0774_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[14\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12191__A2 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12156_ _04813_ _04858_ _04986_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__nor3_2
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06910__A _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6737__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12631__B _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5660_ MuI._1813_ MuI._0246_ MuI._0420_ MuI._1318_ vssd1 vssd1 vccd1 vccd1 MuI._1469_
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11107_ _03809_ _04327_ _03711_ _03857_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._3868__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1534_ AuI._0652_ AuI._0657_ vssd1 vssd1 vccd1 vccd1 AuI._0717_ sky130_fd_sc_hd__and2_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ _04769_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._540_ AuI.pe._393_ AuI.pe._026_ AuI.pe._023_ AuI.pe.significand\[7\] AuI.pe._037_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._098_ sky130_fd_sc_hd__a221o_1
XFILLER_110_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4611_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._0315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5591_ MuI._1377_ MuI._1378_ MuI._1392_ vssd1 vssd1 vccd1 vccd1 MuI._1393_ sky130_fd_sc_hd__and3_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11038_ _06608_ _06546_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__nand2_1
XAuI._1465_ AuI._0646_ AuI._0647_ AuI._0648_ AuI._0649_ AuI._0650_ vssd1 vssd1 vccd1
+ vccd1 AuI._0651_ sky130_fd_sc_hd__o2111ai_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10151__B _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4542_ MuI.b_operand\[21\] MuI._3372_ MuI._0111_ MuI.b_operand\[22\] vssd1 vssd1
+ vccd1 vccd1 MuI._0239_ sky130_fd_sc_hd__a22o_1
XAuI.pe._471_ AuI.pe.significand\[24\] vssd1 vssd1 vccd1 vccd1 AuI.pe._035_ sky130_fd_sc_hd__inv_2
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1396_ net19 net51 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0586_ sky130_fd_sc_hd__mux2_2
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4473_ MuI._0155_ MuI._0160_ MuI._0161_ MuI._0162_ vssd1 vssd1 vccd1 vccd1 MuI._0164_
+ sky130_fd_sc_hd__o31a_1
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _05866_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12359__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6212_ MuI._1274_ MuI._3091_ MuI._1935_ MuI._1932_ vssd1 vssd1 vccd1 vccd1 MuI._2076_
+ sky130_fd_sc_hd__a31o_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3424_ MuI.b_operand\[23\] MuI.b_operand\[26\] MuI._0010_ vssd1 vssd1 vccd1 vccd1
+ MuI._0021_ sky130_fd_sc_hd__and3_1
XFILLER_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11454__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11454__B2 _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6143_ MuI._1998_ MuI._1999_ vssd1 vssd1 vccd1 vccd1 MuI._2001_ sky130_fd_sc_hd__or2b_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1171__A1 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08870__A2 _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6074_ MuI._3067_ MuI._1899_ vssd1 vssd1 vccd1 vccd1 MuI._1925_ sky130_fd_sc_hd__nand2_1
X_07200_ net110 vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__buf_4
XFILLER_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5793__B2 MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12403__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ _00781_ _00797_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__xnor2_2
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4005__B MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5025_ MuI._0765_ MuI._0769_ MuI._0770_ MuI._0653_ vssd1 vssd1 vccd1 vccd1 MuI._0771_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_186_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1517__A AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10229__B_N _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11710__B _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ net112 _03593_ _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__and4_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__B _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07062_ _04004_ _06067_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2_1
XANTENNA__07188__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12822__A _05700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__A_N _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5927_ MuI._1713_ MuI._1762_ MuI._1759_ vssd1 vssd1 vccd1 vccd1 MuI._1763_ sky130_fd_sc_hd__a21o_1
XFILLER_114_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07916__A _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._807_ AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 AuI.pe._346_ sky130_fd_sc_hd__clkinv_2
XANTENNA__12541__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B1 _01988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5858_ MuI._0750_ MuI._1685_ MuI._1686_ vssd1 vssd1 vccd1 vccd1 MuI._1687_ sky130_fd_sc_hd__nand3_1
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07964_ _00275_ _00276_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__nor2_1
XANTENNA__08138__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._738_ AuI.pe._158_ AuI.pe._096_ AuI.pe._119_ AuI.pe._142_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._283_ sky130_fd_sc_hd__a22o_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4809_ MuI._0496_ MuI._0495_ vssd1 vssd1 vccd1 vccd1 MuI._0533_ sky130_fd_sc_hd__and2_1
X_09703_ _02269_ _02316_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__xnor2_2
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08138__B2 _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__A1 _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ _04509_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__buf_6
XMuI._5789_ MuI._0743_ MuI._0742_ MuI._0741_ vssd1 vssd1 vccd1 vccd1 MuI._1611_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07895_ _00511_ _00512_ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__xnor2_1
XAuI.pe._669_ AuI.pe._125_ AuI.pe._384_ AuI.pe._387_ AuI.pe._023_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._218_ sky130_fd_sc_hd__a31o_1
X_09634_ _02272_ _02271_ _06475_ _04111_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__and4bb_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06846_ _03755_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__and3_1
XANTENNA__07361__A2 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09565_ _06491_ _04434_ _04509_ _06492_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22oi_2
X_06777_ _03024_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__and3_1
XANTENNA__13434__A2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11173__A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08466__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _01123_ _01124_ _01131_ _01132_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__nor4_2
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _02120_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__nand3_1
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ _01054_ _01055_ _01062_ _01063_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__or4bb_4
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _00993_ _00994_ _00995_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__or3_1
XFILLER_165_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFuI._082_ FuI.a_operand\[4\] FuI._046_ vssd1 vssd1 vccd1 vccd1 FuI._047_ sky130_fd_sc_hd__and2_1
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07329_ _06599_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__buf_4
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06714__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10340_ _03030_ _03031_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and3_1
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3547__B1 MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _00713_ _00748_ _00746_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__o21ai_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07248__D _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A1 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08377__B2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _04828_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__xor2_2
XFILLER_79_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07826__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06730__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12451__B _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3770__A MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12912_ _05797_ _05798_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__xnor2_1
XAuI._1250_ AuI._0448_ AuI._0451_ vssd1 vssd1 vccd1 vccd1 AuI._0452_ sky130_fd_sc_hd__or2_1
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6264__A2 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07352__A2 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12843_ _05714_ _05715_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__a21oi_1
XAuI._1181_ AuI._0276_ AuI._0385_ AuI._0386_ AuI._0153_ vssd1 vssd1 vccd1 vccd1 AuI._0387_
+ sky130_fd_sc_hd__o211a_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08376__B _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10239__A2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _05648_ _05650_ _05545_ _05611_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o211a_1
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1153__A1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11725_ _04394_ _04393_ _04392_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__a21bo_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09488__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ _02980_ _04972_ _05036_ _00281_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a22o_1
XANTENNA__06905__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ _02884_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__inv_2
XFILLER_128_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _02754_ _02797_ _00385_ _00783_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__and4_1
XFILLER_155_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10183__A_N _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08542__D _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13326_ _06226_ _06176_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10538_ _02229_ _06537_ _00385_ _02431_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a22o_1
XFILLER_155_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0965_ AuI._0171_ AuI._0173_ AuI._0176_ vssd1 vssd1 vccd1 vccd1 AuI._0177_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._6040__B MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__B _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6830_ MuI._2683_ MuI._2701_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI.result\[7\]
+ sky130_fd_sc_hd__nor3b_1
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _06165_ _06122_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__nand2_1
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10469_ _03168_ _03169_ _03158_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07158__D net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0896_ net28 net60 vssd1 vssd1 vccd1 vccd1 AuI._0116_ sky130_fd_sc_hd__nor2_2
XANTENNA_AuI._0895__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6761_ MuI._2588_ MuI._2597_ MuI._2601_ MuI._2679_ vssd1 vssd1 vccd1 vccd1 MuI._2680_
+ sky130_fd_sc_hd__and4_1
XANTENNA__09565__B1 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _05039_ _05040_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a21oi_1
XMuI._3973_ MuI._2971_ MuI._2969_ MuI._2970_ vssd1 vssd1 vccd1 vccd1 MuI._3073_ sky130_fd_sc_hd__nand3_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13188_ _02751_ _06013_ _06014_ _06094_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__a31o_2
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5712_ MuI._2660_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._1526_ sky130_fd_sc_hd__nand2_1
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0967__A1 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6692_ MuI._2383_ MuI._2603_ vssd1 vssd1 vccd1 vccd1 MuI._2604_ sky130_fd_sc_hd__xor2_1
X_12139_ _04967_ _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__nand3_1
XANTENNA__07455__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5643_ MuI._1405_ MuI._1407_ MuI._1402_ vssd1 vssd1 vccd1 vccd1 MuI._1451_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1517_ AuI._0599_ AuI._0692_ vssd1 vssd1 vccd1 vccd1 AuI._0702_ sky130_fd_sc_hd__nand2_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._523_ AuI.pe._020_ AuI.pe._079_ AuI.pe._082_ vssd1 vssd1 vccd1 vccd1 AuI.pe._083_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06700_ _02194_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__buf_6
XFILLER_65_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5574_ MuI._1364_ MuI._1360_ vssd1 vssd1 vccd1 vccd1 MuI._1375_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1448_ AuI._0630_ AuI._0631_ AuI._0623_ AuI._0633_ vssd1 vssd1 vccd1 vccd1 AuI._0634_
+ sky130_fd_sc_hd__or4b_1
X_07680_ _00265_ _00277_ _00297_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__o21ai_4
XAuI.pe._454_ AuI.pe._014_ vssd1 vssd1 vccd1 vccd1 AuI.pe._020_ sky130_fd_sc_hd__clkbuf_4
XMuI._4525_ MuI._0090_ MuI._0214_ vssd1 vssd1 vccd1 vccd1 MuI._0221_ sky130_fd_sc_hd__nor2_1
XFILLER_92_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07471__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1379_ AuI._0552_ AuI._0563_ AuI._0551_ vssd1 vssd1 vccd1 vccd1 AuI._0571_ sky130_fd_sc_hd__and3b_1
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4456_ MuI._0015_ MuI._0139_ MuI._0144_ vssd1 vssd1 vccd1 vccd1 MuI._0145_ sky130_fd_sc_hd__and3_1
X_09350_ _01966_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__nor2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08717__D _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07621__D _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5757__D MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ _00593_ _00595_ _00594_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__o21ai_2
XMuI._4387_ MuI._0064_ MuI._0066_ MuI._0068_ vssd1 vssd1 vccd1 vccd1 MuI._0070_ sky130_fd_sc_hd__and3_1
X_09281_ _06578_ _06579_ _00271_ _04229_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__and4_1
XMuI._6126_ MuI._1883_ MuI._1903_ vssd1 vssd1 vccd1 vccd1 MuI._1982_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._5766__A1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08232_ _06620_ _00445_ _00546_ _00547_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_MuI._5766__B2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06815__A _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3777__B1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6057_ MuI._3125_ MuI._3152_ MuI._1905_ vssd1 vssd1 vccd1 vccd1 MuI._1906_ sky130_fd_sc_hd__a21o_1
X_08163_ _00771_ _00780_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__xnor2_2
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_A net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5008_ MuI._0561_ MuI._0568_ vssd1 vssd1 vccd1 vccd1 MuI._0752_ sky130_fd_sc_hd__xor2_1
XFILLER_162_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6715__A0 MuI._2625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ _05671_ _06414_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__and2_1
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08094_ _00672_ _00711_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__xor2_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07045_ _05906_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__clkbuf_4
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13352__B2 _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11363__B1 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0958__A1 net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08996_ _01365_ _01380_ _01379_ _01372_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a211o_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13104__A1 _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__D _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07947_ _00011_ _00040_ _04789_ _00012_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
XANTENNA__11115__B1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3701__B1 MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07878_ _00493_ _00494_ _00484_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._6246__A2 MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _02233_ _02232_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__xor2_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06829_ net57 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__buf_2
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ _02550_ _04057_ _02178_ _02179_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a31oi_4
XFILLER_197_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11969__A2 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _02100_ _02094_ _02095_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__nand3_1
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _04289_ _04290_ _04088_ _04090_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a211o_1
XFILLER_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ _05344_ _05345_ _05266_ _05236_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a211oi_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06725__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFuI._134_ FuI._018_ net140 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[5\] sky130_fd_sc_hd__dlxtn_1
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12446__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ _04200_ _04201_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11350__B _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13040__B1 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._065_ FuI.a_operand\[25\] net104 FuI.a_operand\[26\] vssd1 vssd1 vccd1 vccd1
+ FuI._033_ sky130_fd_sc_hd__a21o_1
XFILLER_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08598__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__B2 _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__D _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _03902_ _03904_ _04142_ _04143_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__a211oi_4
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13111_ _06011_ _02910_ _04635_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__mux2_1
XFILLER_152_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ _03011_ _03012_ _03008_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a21o_1
XFILLER_152_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4732__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input53_A b_operand[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _05826_ _05910_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2b_1
X_10254_ _02532_ _02559_ _02741_ _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o211a_1
XANTENNA__09474__C _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1071__A0 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10185_ _05209_ _03110_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__and2b_1
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1302_ AuI._0276_ AuI._0390_ AuI._0389_ vssd1 vssd1 vccd1 vccd1 AuI._0500_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1374__A1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1233_ AuI._0435_ AuI._0434_ vssd1 vssd1 vccd1 vccd1 AuI._0436_ sky130_fd_sc_hd__nor2_1
XANTENNA__08752__A1_N _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4310_ MuI._3267_ MuI._3409_ vssd1 vssd1 vccd1 vccd1 MuI._3410_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5290_ MuI._0844_ MuI._1061_ vssd1 vssd1 vccd1 vccd1 MuI._1062_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12826_ _05696_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__xnor2_1
XAuI._1164_ AuI._0271_ AuI._0273_ AuI._0290_ AuI._0291_ AuI._0206_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0371_ sky130_fd_sc_hd__mux4_1
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4241_ MuI._3253_ MuI._3339_ MuI._3338_ MuI._3325_ vssd1 vssd1 vccd1 vccd1 MuI._3341_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_62_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__A1 _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _05631_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nor2_1
XAuI._1095_ AuI._0180_ AuI._0182_ AuI._0185_ AuI._0187_ AuI._0175_ AuI._0205_ vssd1
+ vssd1 vccd1 vccd1 AuI._0305_ sky130_fd_sc_hd__mux4_1
XANTENNA__08825__A2 _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4172_ MuI._2896_ MuI._3271_ vssd1 vssd1 vccd1 vccd1 MuI._3272_ sky130_fd_sc_hd__xor2_1
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _04503_ _04504_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__xor2_1
XFILLER_148_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12688_ _05471_ _05473_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o211ai_4
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11639_ _06434_ _03604_ _06612_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and3_1
XANTENNA__08589__A1 _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08589__B2 _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4971__A2 MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07169__C net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _02833_ _06159_ _02911_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21ba_1
XAuI._0948_ net57 net25 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0160_ sky130_fd_sc_hd__mux2_1
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6813_ MuI._2503_ MuI._2735_ vssd1 vssd1 vccd1 vccd1 MuI.Overflow sky130_fd_sc_hd__nor2_1
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07466__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0879_ net22 net54 vssd1 vssd1 vccd1 vccd1 AuI._0099_ sky130_fd_sc_hd__or2b_1
XMuI._6744_ MuI._2308_ MuI._2475_ vssd1 vssd1 vccd1 vccd1 MuI._2662_ sky130_fd_sc_hd__nor2_1
XFILLER_112_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3956_ MuI._0328_ MuI._2874_ vssd1 vssd1 vccd1 vccd1 MuI._3056_ sky130_fd_sc_hd__and2_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ _01461_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08210__B1 _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07801_ _00416_ _00417_ _00418_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__nand3_1
XFILLER_69_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6675_ MuI._2585_ vssd1 vssd1 vccd1 vccd1 MuI._2586_ sky130_fd_sc_hd__clkinv_2
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3887_ MuI._2983_ MuI._2986_ vssd1 vssd1 vccd1 vccd1 MuI._2987_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08781_ _01397_ _01398_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__and2b_1
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5626_ MuI._1431_ MuI._1413_ MuI._1426_ MuI._1400_ vssd1 vssd1 vccd1 vccd1 MuI._1432_
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07732_ _00344_ _00348_ _00349_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI.pe._541__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._506_ AuI.pe.significand\[4\] AuI.pe._023_ AuI.pe._027_ AuI.pe._062_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._067_ sky130_fd_sc_hd__a22o_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5557_ MuI._1348_ MuI._1349_ MuI._1354_ vssd1 vssd1 vccd1 vccd1 MuI._1356_ sky130_fd_sc_hd__nand3_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07663_ net113 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__buf_4
XFILLER_93_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10320__A1 _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._437_ AuI.pe._003_ vssd1 vssd1 vccd1 vccd1 AuI.pe._004_ sky130_fd_sc_hd__buf_2
XFILLER_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4508_ MuI._0191_ MuI._0195_ MuI._0200_ MuI._0201_ vssd1 vssd1 vccd1 vccd1 MuI._0202_
+ sky130_fd_sc_hd__a211o_1
X_09402_ _01995_ _02017_ _02018_ _02019_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__o211ai_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5488_ MuI._1272_ MuI._1278_ MuI._1279_ vssd1 vssd1 vccd1 vccd1 MuI._1280_ sky130_fd_sc_hd__nor3_1
X_07594_ _06676_ _00025_ _00210_ _00211_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__o211ai_4
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07351__D _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4439_ MuI._0120_ MuI._0125_ vssd1 vssd1 vccd1 vccd1 MuI._0126_ sky130_fd_sc_hd__xnor2_1
X_09333_ _01796_ _01833_ _01834_ _01831_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__o22ai_2
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1668__A2 AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__A _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _01842_ _01810_ _01841_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__nand3_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6109_ MuI._1891_ MuI._1892_ vssd1 vssd1 vccd1 vccd1 MuI._1963_ sky130_fd_sc_hd__nand2_1
XFILLER_178_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08215_ _00824_ _00831_ _00832_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__a21bo_1
X_09195_ _01771_ _01769_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__nor2_1
XFILLER_21_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _00755_ _00762_ _00763_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__nand3_1
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13176__A1_N _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _03378_ _00279_ _04358_ _00083_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__nand4_2
X_07028_ _05724_ _02042_ _05144_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__and3_1
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07807__C _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12813__A2_N _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ _01594_ _01595_ _01596_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10097__B_N _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5675__B1 MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._532__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ _04806_ _04807_ _04675_ _04695_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__o211ai_1
XFILLER_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1356__A1 net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10941_ FuI.Integer\[4\] _06056_ _03674_ _03678_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__D _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10872_ _03602_ _03603_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _05301_ _05306_ _05475_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a211oi_2
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08807__A2 _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1659__A2 AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _05400_ _05401_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__nor2_1
XFILLER_197_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5694__B MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._3495__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11080__B _03828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ _05178_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__or3_4
XFILLER_184_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._117_ FuI._025_ FuI._026_ FuI._028_ vssd1 vssd1 vccd1 vccd1 FuI._029_ sky130_fd_sc_hd__and3_1
XFILLER_200_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12367__A2 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ _04196_ _04198_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__nand3_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10378__A1 _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12904__B _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _04124_ _04121_ _04123_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nand3_2
XANTENNA__10705__A _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12119__A2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ _00698_ _00702_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a211oi_1
XFILLER_180_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08820__D net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ _03913_ _03910_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3810_ MuI._2908_ MuI._2909_ vssd1 vssd1 vccd1 vccd1 MuI._2910_ sky130_fd_sc_hd__and2b_1
XFILLER_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12342__D _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ _05746_ _05835_ _05836_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a21oi_1
XMuI._4790_ MuI._0458_ MuI._0461_ vssd1 vssd1 vccd1 vccd1 MuI._0512_ sky130_fd_sc_hd__and2_1
X_10237_ _02824_ _02919_ _02920_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__o211a_1
XMuI._3741_ MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 MuI._2841_ sky130_fd_sc_hd__clkbuf_4
XFILLER_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10168_ _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__inv_2
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6460_ MuI._2343_ MuI._2345_ MuI._2348_ vssd1 vssd1 vccd1 vccd1 MuI._2349_ sky130_fd_sc_hd__o21ai_1
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3672_ MuI._2462_ MuI._2561_ MuI._2506_ vssd1 vssd1 vccd1 vccd1 MuI._2743_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._523__A2 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10099_ _02771_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__and2_1
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5411_ MuI._3362_ MuI._3262_ MuI._0020_ MuI._0085_ vssd1 vssd1 vccd1 vccd1 MuI._1195_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1347__A1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6391_ MuI._2271_ MuI._1975_ MuI._2272_ vssd1 vssd1 vccd1 vccd1 MuI._2273_ sky130_fd_sc_hd__a21o_1
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6046__A MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3692__A2 MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5342_ MuI._1084_ MuI._1118_ vssd1 vssd1 vccd1 vccd1 MuI._1119_ sky130_fd_sc_hd__xnor2_1
XAuI._1216_ AuI._0419_ vssd1 vssd1 vccd1 vccd1 AuI._0420_ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5273_ MuI._1037_ MuI._1041_ MuI._1042_ vssd1 vssd1 vccd1 vccd1 MuI._1044_ sky130_fd_sc_hd__nand3_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _03271_ _00153_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__and2_1
XAuI._1147_ AuI._0189_ AuI._0236_ AuI._0198_ AuI._0202_ AuI._0307_ vssd1 vssd1 vccd1
+ vccd1 AuI._0355_ sky130_fd_sc_hd__a311o_1
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4224_ MuI._3209_ MuI._3323_ vssd1 vssd1 vccd1 vccd1 MuI._3324_ sky130_fd_sc_hd__or2_1
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1078_ AuI._0263_ AuI._0275_ AuI._0287_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0289_
+ sky130_fd_sc_hd__a211o_1
XFILLER_188_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09379__C net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4155_ MuI._3215_ MuI._3254_ vssd1 vssd1 vccd1 vccd1 MuI._3255_ sky130_fd_sc_hd__xor2_1
X_08000_ _00615_ _00614_ _00616_ _00617_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__nand4_2
XMuI._4086_ MuI.a_operand\[22\] MuI._2894_ MuI._2892_ MuI._3185_ vssd1 vssd1 vccd1
+ vccd1 MuI._3186_ sky130_fd_sc_hd__and4_1
XFILLER_129_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1525__A AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13307__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09951_ _02341_ _02340_ _02603_ _02610_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__nand4_1
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ _06620_ _04456_ _01351_ _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a31o_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4988_ MuI._0727_ MuI._0729_ vssd1 vssd1 vccd1 vccd1 MuI._0730_ sky130_fd_sc_hd__and2_1
X_09882_ _02537_ _02531_ _02535_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__nor3_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A1 _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11869__B2 _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6727_ MuI._2642_ vssd1 vssd1 vccd1 vccd1 MuI._2643_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__08734__A1 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3939_ MuI._3038_ vssd1 vssd1 vccd1 vccd1 MuI._3039_ sky130_fd_sc_hd__inv_2
X_08833_ _01332_ _02334_ _06604_ _06580_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__and4_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10541__A1 _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6658_ MuI._0999_ MuI._2482_ MuI._2483_ MuI._2566_ vssd1 vssd1 vccd1 vccd1 MuI._2567_
+ sky130_fd_sc_hd__or4_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _01374_ _01376_ _01375_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12818__B1 _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5609_ MuI._1412_ vssd1 vssd1 vccd1 vccd1 MuI._1413_ sky130_fd_sc_hd__inv_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _00331_ _00330_ _00329_ _00328_ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__o211a_1
XMuI._6589_ MuI.b_operand\[23\] MuI._2488_ MuI._2489_ MuI._2490_ vssd1 vssd1 vccd1
+ vccd1 MuI._2491_ sky130_fd_sc_hd__a31o_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11097__A2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _01214_ _01274_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07646_ _00091_ _00263_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__nor2_1
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6082__B1 MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._817__A3 AuI.pe._070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13243__B1 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07577_ _00192_ _00193_ _00194_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__nand3_1
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09316_ _01931_ _01932_ _01933_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__o21bai_1
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _01855_ _01856_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__or4_4
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4396__B1 MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09178_ _01789_ _01794_ _01784_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a211oi_2
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _00744_ _00745_ _00430_ _00433_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__o211ai_1
XANTENNA__11021__A2 _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ _03881_ _03891_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__and3_2
XFILLER_162_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1026__A0 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 ALU_Output[18] sky130_fd_sc_hd__buf_2
X_11071_ _03740_ _03818_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__xnor2_2
XANTENNA_MuI._3481__C MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 ALU_Output[28] sky130_fd_sc_hd__buf_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08725__A1 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10022_ _02685_ _02690_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08725__B2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5112__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A2_N _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A a_operand[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _04786_ _04787_ _04788_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._680__B AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10924_ _03294_ _03485_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nor2_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08665__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1001_ AuI._0153_ AuI._0210_ AuI._0212_ vssd1 vssd1 vccd1 vccd1 AuI._0213_ sky130_fd_sc_hd__a21o_1
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _03582_ _03583_ _03584_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a21o_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__B_N _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10786_ _03375_ _03338_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or2b_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _05381_ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__nand2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nand2_1
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06913__A _04489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5960_ MuI._0765_ MuI._0766_ vssd1 vssd1 vccd1 vccd1 MuI._1799_ sky130_fd_sc_hd__and2b_1
XFILLER_126_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _03809_ _04467_ _04110_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and3_1
XANTENNA__08413__B1 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ _05232_ _05233_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__and3_1
XFILLER_181_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4911_ MuI._0635_ MuI._0644_ vssd1 vssd1 vccd1 vccd1 MuI._0645_ sky130_fd_sc_hd__xnor2_1
XANTENNA_output84_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5891_ MuI._0719_ MuI._0721_ vssd1 vssd1 vccd1 vccd1 MuI._1723_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__xnor2_4
XFILLER_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10771__A1 _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._771_ AuI.pe._314_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[22\] sky130_fd_sc_hd__clkbuf_1
XMuI._4842_ MuI._0561_ MuI._0568_ vssd1 vssd1 vccd1 vccd1 MuI._0569_ sky130_fd_sc_hd__and2_1
XANTENNA_AuI._1017__A0 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11269_ _02840_ _05585_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__nand2_1
XANTENNA__08716__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13008_ _05800_ _05802_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__o21a_1
XMuI._4773_ MuI._0325_ MuI._0492_ vssd1 vssd1 vccd1 vccd1 MuI._0494_ sky130_fd_sc_hd__or2_1
XFILLER_95_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07744__A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13465__B _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6512_ MuI._2000_ MuI._2099_ MuI._1989_ vssd1 vssd1 vccd1 vccd1 MuI._2406_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3724_ MuI._2819_ MuI._2823_ vssd1 vssd1 vccd1 vccd1 MuI._2824_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10170__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09381__D _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6443_ MuI._2320_ MuI._2328_ MuI._2295_ MuI._2329_ vssd1 vssd1 vccd1 vccd1 MuI._2331_
+ sky130_fd_sc_hd__a211oi_2
XMuI._3655_ MuI._2517_ MuI._2528_ MuI._2539_ MuI._2550_ vssd1 vssd1 vccd1 vccd1 MuI._2561_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07500_ _00115_ _00116_ _00117_ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__and3_1
XFILLER_208_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6374_ MuI._2090_ MuI._2254_ vssd1 vssd1 vccd1 vccd1 MuI._2255_ sky130_fd_sc_hd__nor2_1
XFILLER_208_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3586_ MuI._1791_ vssd1 vssd1 vccd1 vccd1 MuI._1802_ sky130_fd_sc_hd__buf_2
XANTENNA__10117__A_N _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _00920_ _01097_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5325_ MuI._1085_ MuI._1086_ MuI._1100_ vssd1 vssd1 vccd1 vccd1 MuI._1101_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4008__B MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12809__B _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07431_ net43 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__buf_6
XFILLER_196_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4614__A1 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12097__A _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5256_ MuI._1022_ MuI._1023_ MuI._1017_ vssd1 vssd1 vccd1 vccd1 MuI._1025_ sky130_fd_sc_hd__a21o_1
X_07362_ net106 vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__buf_4
XFILLER_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3847__B MuI._0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4207_ MuI.b_operand\[3\] vssd1 vssd1 vccd1 vccd1 MuI._3307_ sky130_fd_sc_hd__buf_2
X_09101_ _01713_ _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__and2_1
XMuI._5187_ MuI._0819_ MuI._0822_ MuI._0824_ MuI._0826_ vssd1 vssd1 vccd1 vccd1 MuI._0949_
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11251__A2 _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07293_ _06593_ _04972_ _06589_ _06590_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4138_ MuI._1153_ MuI._2363_ MuI._2385_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._3238_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _01647_ _01648_ _01649_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a21o_1
XANTENNA__07919__A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08741__C _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4069_ MuI._2865_ MuI._2924_ vssd1 vssd1 vccd1 vccd1 MuI._3169_ sky130_fd_sc_hd__xor2_2
XANTENNA__11003__A2 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07758__A2 _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1405__D AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4397__C MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1008__A0 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ _02585_ _02595_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI.pe._735__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07654__A _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09865_ _02484_ _02486_ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a21o_1
XANTENNA_input8_A a_operand[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__A1 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _01408_ _01431_ _01432_ _01433_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nand4_2
XANTENNA__09380__B2 _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _02444_ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__or2_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ _01342_ _01347_ _01364_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__a21o_2
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6117__C MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08678_ _00986_ _00987_ _01002_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__a21oi_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07629_ _00228_ _00229_ _00246_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__and3_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10640_ _03353_ _03354_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__xnor2_4
XFILLER_198_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08635__D _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07446__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__A3 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _03106_ _03104_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__and2b_1
XANTENNA__07446__B2 _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _05039_ _05151_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__o21a_1
XANTENNA__07829__A _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13290_ _06066_ _06070_ _06139_ _06062_ _06061_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a2111o_1
XFILLER_155_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06733__A _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3773__A MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ _06444_ _06442_ _00534_ _06525_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and4_1
XFILLER_135_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10255__A _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3592__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3592__B2 MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08370__D net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _02848_ _05003_ _04161_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__o21a_1
XFILLER_123_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11123_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__and2_1
XFILLER_150_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1550_ AuI._0606_ AuI._0729_ AuI._0730_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[5\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4100__C MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _06565_ _03082_ _00789_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__and3_1
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1481_ AuI._0635_ AuI._0637_ vssd1 vssd1 vccd1 vccd1 AuI._0667_ sky130_fd_sc_hd__and2b_1
XFILLER_77_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10005_ _02670_ _02668_ _02667_ _01866_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09371__B2 _01988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__C _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12258__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3440_ MuI.a_operand\[27\] MuI.b_operand\[27\] vssd1 vssd1 vccd1 vccd1 MuI._0196_
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__A _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _00058_ _03449_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nand2_1
XANTENNA__07134__B1 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06908__A _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08826__C net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ _03641_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nor2_1
X_11887_ _04525_ _04546_ _04696_ _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a211o_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__B1 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5110_ MuI._0857_ MuI._0851_ MuI._0852_ vssd1 vssd1 vccd1 vccd1 MuI._0864_ sky130_fd_sc_hd__nand3_1
XFILLER_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6090_ MuI._0867_ MuI._2594_ vssd1 vssd1 vccd1 vccd1 MuI._1942_ sky130_fd_sc_hd__nand2_1
X_10838_ _03565_ _03566_ _03567_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21o_1
XFILLER_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5041_ MuI._0015_ MuI._0139_ MuI._0144_ vssd1 vssd1 vccd1 vccd1 MuI._0788_ sky130_fd_sc_hd__nand3_1
XFILLER_60_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ _02129_ _03306_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__nor2_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07988__A2 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ FuI.Integer\[16\] _02931_ _02719_ _05058_ _05365_ vssd1 vssd1 vccd1 vccd1
+ _05366_ sky130_fd_sc_hd__a221o_1
X_13488_ _02812_ _06354_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__and2_1
XFILLER_139_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12439_ _00676_ _06568_ _03047_ _00506_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10165__A _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12194__B1 _00555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__C _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5943_ MuI._1777_ MuI._1778_ MuI._1773_ MuI._1774_ vssd1 vssd1 vccd1 vccd1 MuI._1781_
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._823_ AuI.pe._339_ AuI.pe._344_ AuI.pe._357_ vssd1 vssd1 vccd1 vccd1 AuI.pe._361_
+ sky130_fd_sc_hd__o21a_1
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11941__B1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5874_ MuI._1667_ MuI._1702_ MuI._1704_ vssd1 vssd1 vccd1 vccd1 MuI._1705_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI.pe._585__B AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout109 net63 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_6
X_07980_ _00260_ _00591_ _00597_ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._754_ AuI.pe.significand\[8\] AuI.pe._375_ AuI.pe._297_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._298_ sky130_fd_sc_hd__or3_1
XMuI._4825_ MuI._0549_ MuI._0550_ vssd1 vssd1 vccd1 vccd1 MuI._0551_ sky130_fd_sc_hd__and2_1
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06931_ _04682_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._685_ AuI.pe._142_ AuI.pe._086_ AuI.pe._232_ vssd1 vssd1 vccd1 vccd1 AuI.pe._233_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5403__A MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4756_ MuI._0340_ MuI._0474_ vssd1 vssd1 vccd1 vccd1 MuI._0475_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4945__C MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _02251_ _02242_ _02250_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__nand3_1
XFILLER_110_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06862_ _03939_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[0\] sky130_fd_sc_hd__clkbuf_2
XANTENNA__11427__C _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3707_ MuI._2780_ MuI._2805_ MuI._2795_ vssd1 vssd1 vccd1 vccd1 MuI._2807_ sky130_fd_sc_hd__nand3_1
X_08601_ _00988_ _00990_ _00989_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4687_ MuI._0341_ MuI._0363_ vssd1 vssd1 vccd1 vccd1 MuI._0399_ sky130_fd_sc_hd__xor2_1
X_09581_ _02143_ _02188_ _02211_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a211o_1
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06793_ _03196_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[20\] sky130_fd_sc_hd__clkbuf_2
XFILLER_209_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6426_ MuI._2250_ MuI._2252_ MuI._2266_ vssd1 vssd1 vccd1 vccd1 MuI._2312_ sky130_fd_sc_hd__o21ai_1
XMuI._3638_ MuI.a_operand\[7\] vssd1 vssd1 vccd1 vccd1 MuI._2374_ sky130_fd_sc_hd__clkbuf_4
X_08532_ _01144_ _01149_ _03400_ _03906_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__o211a_1
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6357_ MuI._2234_ MuI._2202_ MuI._2191_ vssd1 vssd1 vccd1 vccd1 MuI._2236_ sky130_fd_sc_hd__nor3_1
XANTENNA__08736__C _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3569_ MuI._0856_ MuI._1604_ vssd1 vssd1 vccd1 vccd1 MuI._1615_ sky130_fd_sc_hd__xnor2_2
X_08463_ _01079_ _01080_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__nor2_1
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5308_ MuI._1073_ MuI._1079_ MuI._1080_ vssd1 vssd1 vccd1 vccd1 MuI._1082_ sky130_fd_sc_hd__nor3_1
XFILLER_168_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ net8 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6288_ MuI._2158_ MuI._2159_ vssd1 vssd1 vccd1 vccd1 MuI._2160_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _00840_ _01011_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._653__A1 AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5239_ MuI._1004_ MuI._1005_ vssd1 vssd1 vccd1 vccd1 MuI._1006_ sky130_fd_sc_hd__and2b_1
X_07345_ _06643_ _06644_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__or3_1
XANTENNA__09848__B _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07649__A _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5792__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _06575_ _06574_ _06533_ _06511_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__o211ai_2
XFILLER_192_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _01555_ _01554_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__and2b_1
XFILLER_191_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07600__A1 _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07600__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07384__A _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _02394_ _02443_ _02347_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12488__A1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3877__A2 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__B _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08199__B _00664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12440__D _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5079__A1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _02302_ _02345_ net115 _06436_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__and4_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5079__B2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07364__B1 _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _02388_ _03971_ _02410_ _02427_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a31o_1
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07831__B _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ _04310_ _04484_ _04486_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a21o_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12790_ _05667_ _05668_ _06427_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06728__A _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _04537_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a21oi_1
XFILLER_82_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4590__C MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11672_ _04464_ _04465_ _04446_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10623_ _03157_ _03177_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a21boi_2
X_13411_ _06286_ _06324_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11215__A2 _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3801__A2 MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07559__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ _06252_ _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__and2b_1
XFILLER_183_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12963__A2 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ _00791_ _03090_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__o21a_1
XAuI._0981_ AuI._0155_ AuI._0158_ AuI._0160_ AuI._0166_ vssd1 vssd1 vccd1 vccd1 AuI._0193_
+ sky130_fd_sc_hd__or4_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13273_ _03809_ _05713_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__nand2_1
XFILLER_155_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ _03182_ _03187_ _03188_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__nand3_1
XFILLER_108_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12176__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12715__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ _05057_ _05059_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nand3b_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10726__A1 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10726__B2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1602_ AuI.pe.Significand\[14\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0774_
+ sky130_fd_sc_hd__or2_1
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _04813_ _04858_ _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o21a_2
XANTENNA_AuI._0864__A2_N net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _03708_ _03710_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__and2b_1
XAuI._1533_ AuI._0713_ vssd1 vssd1 vccd1 vccd1 AuI._0716_ sky130_fd_sc_hd__inv_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12086_ _04910_ _04911_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._3868__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4610_ MuI._0312_ MuI._0313_ vssd1 vssd1 vccd1 vccd1 MuI._0314_ sky130_fd_sc_hd__nor2_1
XMuI._5590_ MuI._1382_ MuI._1390_ MuI._1391_ vssd1 vssd1 vccd1 vccd1 MuI._1392_ sky130_fd_sc_hd__a21o_1
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11037_ _03781_ _03782_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__nor2_1
XFILLER_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1464_ AuI._0392_ AuI._0395_ vssd1 vssd1 vccd1 vccd1 AuI._0650_ sky130_fd_sc_hd__xnor2_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._470_ AuI.pe._028_ AuI.pe._023_ AuI.pe._027_ AuI.pe._033_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._034_ sky130_fd_sc_hd__a22o_1
XMuI._4541_ MuI._0236_ MuI._0237_ vssd1 vssd1 vccd1 vccd1 MuI._0238_ sky130_fd_sc_hd__nor2_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1395_ AuI._0576_ AuI._0583_ vssd1 vssd1 vccd1 vccd1 AuI._0585_ sky130_fd_sc_hd__or2_1
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4472_ MuI._0151_ MuI._0154_ vssd1 vssd1 vccd1 vccd1 MuI._0162_ sky130_fd_sc_hd__nand2_1
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6211_ MuI._2034_ MuI._2040_ MuI._2039_ vssd1 vssd1 vccd1 vccd1 MuI._2075_ sky130_fd_sc_hd__a21o_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ _05877_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__xor2_1
XMuI._3423_ MuI.b_operand\[28\] MuI.b_operand\[27\] MuI.b_operand\[30\] MuI.b_operand\[29\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0010_ sky130_fd_sc_hd__and4_1
XANTENNA__12359__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3678__A MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11454__A2 _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _04654_ _04602_ _04753_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a211oi_4
XFILLER_33_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6142_ MuI._1911_ MuI._1914_ vssd1 vssd1 vccd1 vccd1 MuI._1999_ sky130_fd_sc_hd__xnor2_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6073_ MuI._1921_ MuI._1922_ vssd1 vssd1 vccd1 vccd1 MuI._1924_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__A1 _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5793__A2 MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__B2 _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5024_ MuI._0613_ MuI._0615_ MuI._0651_ MuI._0652_ vssd1 vssd1 vccd1 vccd1 MuI._0770_
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4005__C MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07130_ net126 vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08083__A1 _00698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07830__A1 _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4302__A MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5926_ MuI._1646_ MuI._1711_ vssd1 vssd1 vccd1 vccd1 MuI._1762_ sky130_fd_sc_hd__or2_1
XFILLER_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11719__A _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._806_ AuI.pe._391_ vssd1 vssd1 vccd1 vccd1 AuI.pe._345_ sky130_fd_sc_hd__inv_2
XFILLER_102_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12541__C _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5857_ MuI._0747_ MuI._0748_ MuI._0749_ vssd1 vssd1 vccd1 vccd1 MuI._1686_ sky130_fd_sc_hd__a21o_1
XFILLER_101_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _00570_ _00577_ _00578_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__and3_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._737_ AuI.pe._170_ AuI.pe._399_ AuI.pe._281_ AuI.pe.significand\[20\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._282_ sky130_fd_sc_hd__a22o_1
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4808_ MuI._0529_ MuI._0531_ vssd1 vssd1 vccd1 vccd1 MuI._0532_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08138__A2 _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09702_ _02340_ _02344_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__xnor2_1
X_06914_ net36 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__buf_4
XANTENNA__13131__A2 _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5788_ MuI._1526_ MuI._1529_ MuI._1528_ vssd1 vssd1 vccd1 vccd1 MuI._1610_ sky130_fd_sc_hd__o21bai_1
XANTENNA_AuI.pe._571__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07894_ _06432_ _06438_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__nor2_1
XFILLER_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._668_ AuI.pe._072_ AuI.pe._133_ AuI.pe._173_ AuI.pe._045_ AuI.pe._216_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._217_ sky130_fd_sc_hd__a221o_1
XFILLER_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4739_ MuI._0439_ MuI._0455_ vssd1 vssd1 vccd1 vccd1 MuI._0456_ sky130_fd_sc_hd__or2_1
XFILLER_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07932__A _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ _02151_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__clkbuf_2
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _00162_ _00287_ _00267_ _00164_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22oi_2
XANTENNA__11693__A2 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._599_ AuI.pe._105_ AuI.pe._004_ AuI.pe._022_ AuI.pe._378_ AuI.pe._152_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._153_ sky130_fd_sc_hd__a221o_1
XFILLER_209_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _06488_ _00072_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__nand2_1
XFILLER_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06776_ _03013_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__buf_6
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6409_ MuI._2291_ MuI._2292_ vssd1 vssd1 vccd1 vccd1 MuI._2293_ sky130_fd_sc_hd__xor2_1
XFILLER_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ _01123_ _01124_ _01131_ _01132_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__o22a_1
XANTENNA_MuI._3588__A MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__B _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08446_ _01054_ _01055_ _01062_ _01063_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._626__A1 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._150_ FuI._013_ net156 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[21\] sky130_fd_sc_hd__dlxtn_1
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4488__B_N MuI._0166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _06515_ net133 _06581_ _06519_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a22oi_2
XFILLER_196_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._081_ FuI._035_ FuI._043_ FuI._045_ vssd1 vssd1 vccd1 vccd1 FuI._046_ sky130_fd_sc_hd__or3_1
XFILLER_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07379__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07328_ net121 _04843_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nand2_4
XFILLER_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07259_ net106 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__buf_6
XFILLER_192_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3547__A1 MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3547__B2 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ _00691_ _02955_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a21boi_4
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12732__B _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3770__B MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11348__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11133__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ _05696_ _05705_ _05704_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a21boi_1
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12881__A1 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12881__B2 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__xor2_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1180_ AuI._0236_ AuI._0315_ AuI._0208_ vssd1 vssd1 vccd1 vccd1 AuI._0386_ sky130_fd_sc_hd__a21o_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3498__A MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05545_ _05611_ _05648_ _05650_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a211oi_2
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11724_ _04521_ _04518_ _04519_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__nand3_1
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _04202_ _04205_ _04203_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__o21bai_1
XFILLER_30_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09488__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10708__A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10606_ _03317_ _02883_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or2_1
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11586_ _00878_ _05767_ _03257_ _00877_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__a22oi_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10537_ _03081_ _03084_ _03083_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a21bo_1
X_13325_ _06234_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__or2_1
XAuI._0964_ AuI._0175_ vssd1 vssd1 vccd1 vccd1 AuI._0176_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12923__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10468_ _03158_ _03168_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__and3_1
X_13256_ _06118_ _06120_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or2b_1
XFILLER_136_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06921__A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0895_ net28 net60 vssd1 vssd1 vccd1 vccd1 AuI._0115_ sky130_fd_sc_hd__and2_1
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6760_ MuI._2621_ MuI._2626_ vssd1 vssd1 vccd1 vccd1 MuI._2679_ sky130_fd_sc_hd__and2_1
XANTENNA__09565__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3972_ MuI._2967_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._3072_ sky130_fd_sc_hd__and2_1
XANTENNA__09565__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12207_ _00217_ _05948_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__and3_1
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _03134_ _06072_ _06073_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__a31o_1
X_10399_ _00795_ _00796_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__or2b_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5711_ MuI._1038_ MuI._1040_ MuI._1039_ vssd1 vssd1 vccd1 vccd1 MuI._1525_ sky130_fd_sc_hd__o21bai_1
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6691_ MuI._1996_ MuI._2602_ MuI._2394_ vssd1 vssd1 vccd1 vccd1 MuI._2603_ sky130_fd_sc_hd__a21oi_2
X_12138_ _04965_ _04966_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__a21o_1
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__C _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5642_ MuI._1334_ MuI._1448_ vssd1 vssd1 vccd1 vccd1 MuI._1449_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1516_ AuI._0692_ vssd1 vssd1 vccd1 vccd1 AuI._0701_ sky130_fd_sc_hd__buf_2
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12069_ _02844_ _04893_ _02713_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._522_ AuI.pe._028_ AuI.pe._066_ AuI.pe._054_ AuI.pe._055_ AuI.pe._081_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._082_ sky130_fd_sc_hd__a221o_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5573_ MuI._1368_ MuI._1369_ MuI._1365_ MuI._1367_ vssd1 vssd1 vccd1 vccd1 MuI._1374_
+ sky130_fd_sc_hd__a211o_1
XAuI._1447_ AuI._0624_ AuI._0632_ vssd1 vssd1 vccd1 vccd1 AuI._0633_ sky130_fd_sc_hd__nor2_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._453_ AuI.exp_a AuI.pe._019_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[0\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4524_ MuI._0216_ MuI._0219_ vssd1 vssd1 vccd1 vccd1 MuI._0220_ sky130_fd_sc_hd__or2_1
XFILLER_93_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1378_ AuI._0528_ AuI._0545_ AuI._0551_ AuI._0563_ vssd1 vssd1 vccd1 vccd1 AuI._0570_
+ sky130_fd_sc_hd__and4_1
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4455_ MuI._0140_ MuI._0143_ vssd1 vssd1 vccd1 vccd1 MuI._0144_ sky130_fd_sc_hd__or2b_1
XFILLER_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08300_ _00916_ _00917_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4386_ MuI._0064_ MuI._0066_ MuI._0068_ vssd1 vssd1 vccd1 vccd1 MuI._0069_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09280_ _01794_ _01896_ _01897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__nand3_1
XFILLER_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6125_ MuI._1962_ MuI._1980_ vssd1 vssd1 vccd1 vccd1 MuI._1981_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4016__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._608__B2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08231_ _00835_ _00846_ _00847_ _00848_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__a211oi_4
XFILLER_166_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5766__A2 MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08935__A1_N _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3777__A1 MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6056_ MuI._3149_ MuI._3151_ vssd1 vssd1 vccd1 vccd1 MuI._1905_ sky130_fd_sc_hd__nor2_1
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3777__B2 MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ _00778_ _00779_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__and2b_1
XANTENNA__07199__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5007_ MuI._0747_ MuI._0750_ vssd1 vssd1 vccd1 vccd1 MuI._0751_ sky130_fd_sc_hd__nand2_1
XANTENNA__10938__A1 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07113_ _06420_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[25\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10938__B2 _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6715__A1 MuI._2629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08093_ _00673_ _00710_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__xnor2_2
XFILLER_162_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout116_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07044_ _05895_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__clkbuf_4
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13352__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__A _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10353__A _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5909_ MuI._0685_ MuI._1690_ MuI._1691_ vssd1 vssd1 vccd1 vccd1 MuI._1743_ sky130_fd_sc_hd__or3_1
XFILLER_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ _01609_ _01610_ _01605_ _01608_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__o211a_1
XANTENNA__13104__A2 _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07946_ _00545_ _00561_ _00562_ _00563_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a211oi_4
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3701__B2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07662__A _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _00484_ _00493_ _00494_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__and3_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09616_ _02238_ _02239_ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__and3_1
X_06828_ _03572_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[27\] sky130_fd_sc_hd__clkbuf_1
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ _06564_ _02474_ _04100_ _04165_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__and4_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06759_ net121 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__buf_6
XFILLER_197_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09478_ _02045_ _02102_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__nor2_1
XANTENNA__08493__A _00918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08429_ _01043_ _01045_ _01044_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a21o_1
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0894__A1 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFuI._133_ FuI._017_ net139 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[4\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ _04206_ _04216_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13040__B2 _05926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08598__A2 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _04140_ _04141_ _03989_ _03991_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__o211a_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _02780_ _05993_ _02783_ _05859_ _02781_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__o221ai_1
X_10322_ _03008_ _03011_ _03012_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__nand3_1
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06741__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ _02751_ _05861_ _05862_ _05937_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__a31o_4
X_10253_ _02216_ _03928_ _04004_ _02118_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__a22o_1
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09474__D _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__B1 _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A b_operand[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _02863_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__nor2_2
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1071__A1 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1323__D AuI._0519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5142__B1 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1301_ AuI._0438_ AuI._0383_ vssd1 vssd1 vccd1 vccd1 AuI._0499_ sky130_fd_sc_hd__nor2_1
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1232_ AuI._0427_ AuI._0428_ vssd1 vssd1 vccd1 vccd1 AuI._0435_ sky130_fd_sc_hd__and2b_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nand2_1
XAuI._1163_ AuI._0330_ AuI._0281_ AuI._0369_ AuI._0153_ vssd1 vssd1 vccd1 vccd1 AuI._0370_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4240_ MuI._3325_ MuI._3338_ MuI._3339_ MuI._3253_ vssd1 vssd1 vccd1 vccd1 MuI._3340_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12082__A2 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _03539_ _00678_ _06666_ _00398_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__and4_1
XAuI._1094_ AuI._0261_ AuI._0289_ AuI._0296_ AuI._0213_ AuI._0250_ vssd1 vssd1 vccd1
+ vccd1 AuI._0304_ sky130_fd_sc_hd__a32o_1
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4171_ MuI._2883_ MuI._2887_ MuI._2891_ MuI._2893_ vssd1 vssd1 vccd1 vccd1 MuI._3271_
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3956__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11707_ _02851_ _05777_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__nand2_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10438__A _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _05555_ _05556_ _05492_ _05466_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._4956__B1 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ _04045_ _04048_ _04218_ _04219_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a211o_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08589__A2 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _04352_ _04353_ _04354_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or3_1
XANTENNA__07169__D _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12790__B1 _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13308_ _02833_ _06158_ _02913_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__o21a_1
XAuI._0947_ AuI._0158_ AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 AuI._0159_ sky130_fd_sc_hd__or2b_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6812_ MuI._2504_ MuI._2735_ vssd1 vssd1 vccd1 vccd1 MuI.Underflow sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._3691__A MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _05671_ _02719_ _02722_ _03454_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__a221o_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0878_ net54 net22 vssd1 vssd1 vccd1 vccd1 AuI._0098_ sky130_fd_sc_hd__or2b_1
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6743_ MuI._2657_ MuI._2659_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2661_ sky130_fd_sc_hd__mux2_1
XFILLER_124_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3955_ MuI._0581_ MuI._2898_ vssd1 vssd1 vccd1 vccd1 MuI._3055_ sky130_fd_sc_hd__nand2_1
XANTENNA__08210__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08210__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11896__A2 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5133__B1 MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6674_ MuI._2582_ MuI._2584_ vssd1 vssd1 vccd1 vccd1 MuI._2585_ sky130_fd_sc_hd__or2b_1
XANTENNA_AuI.pe._593__B AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _00189_ _00190_ _00191_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__o21bai_1
XMuI._3886_ MuI._2984_ MuI._2985_ vssd1 vssd1 vccd1 vccd1 MuI._2986_ sky130_fd_sc_hd__nor2_1
X_08780_ _00029_ _00271_ _04229_ _00028_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a22o_1
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5625_ MuI._1400_ MuI._1410_ vssd1 vssd1 vccd1 vccd1 MuI._1431_ sky130_fd_sc_hd__nor2_1
XFILLER_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__A2_N _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _03486_ _04186_ _00346_ _00347_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a22o_1
XAuI.pe._505_ AuI.pe._002_ vssd1 vssd1 vccd1 vccd1 AuI.pe._066_ sky130_fd_sc_hd__buf_2
XFILLER_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5556_ MuI._1348_ MuI._1349_ MuI._1354_ vssd1 vssd1 vccd1 vccd1 MuI._1355_ sky130_fd_sc_hd__a21o_1
XFILLER_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ _00278_ _00279_ _04035_ _06433_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__and4_1
XAuI.pe._436_ AuI.pe._000_ AuI.pe._368_ vssd1 vssd1 vccd1 vccd1 AuI.pe._003_ sky130_fd_sc_hd__nor2_1
XFILLER_92_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4507_ MuI._0176_ MuI._0197_ MuI._0199_ vssd1 vssd1 vccd1 vccd1 MuI._0201_ sky130_fd_sc_hd__and3_1
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10320__A2 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09401_ _01946_ _01948_ _01949_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__or3_1
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5487_ MuI._1270_ MuI._1271_ MuI._1260_ MuI._1269_ vssd1 vssd1 vccd1 vccd1 MuI._1279_
+ sky130_fd_sc_hd__o211a_1
X_07593_ _00186_ _00187_ _00209_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__or3_1
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4438_ MuI._0123_ MuI._0124_ vssd1 vssd1 vccd1 vccd1 MuI._0125_ sky130_fd_sc_hd__nor2_1
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09332_ _01946_ _01948_ _01949_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__nor3_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06826__A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4369_ MuI._3393_ MuI._3411_ vssd1 vssd1 vccd1 vccd1 MuI._0050_ sky130_fd_sc_hd__xor2_2
XANTENNA_MuI._3866__A MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _01850_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__xor2_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6242__A MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6108_ MuI._1958_ MuI._1961_ vssd1 vssd1 vccd1 vccd1 MuI._1962_ sky130_fd_sc_hd__xnor2_1
X_08214_ _00825_ _00830_ _00826_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__nand3_1
XFILLER_119_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _01693_ _01685_ _01692_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__nand3_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6039_ MuI._0581_ MuI._2851_ vssd1 vssd1 vccd1 vccd1 MuI._1886_ sky130_fd_sc_hd__nand2_1
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _00759_ _00760_ _00761_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__a21o_1
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._144__150 vssd1 vssd1 vccd1 vccd1 FuI._144__150/HI net150 sky130_fd_sc_hd__conb_1
X_08076_ _03432_ _04358_ _00083_ _00278_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__a22o_1
XFILLER_134_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ _05713_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10083__A _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07807__D _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11907__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5675__A1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08978_ _06494_ _06495_ net11 net133 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and4_1
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5675__B2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07392__A _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1440__B AuI._0506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ _02658_ _04896_ _04961_ _02593_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a22oi_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _04262_ _03675_ _02721_ _02345_ _03677_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a221o_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ net121 _06477_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nand2_1
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ _05473_ _05474_ _05335_ _05398_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__o211a_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12064__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06736__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3776__A MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ _00299_ _00231_ _06537_ _00385_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__and4_1
XFILLER_185_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0867__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _05324_ _05325_ _05308_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a21oi_1
XFuI._116_ FuI._053_ FuI._027_ vssd1 vssd1 vccd1 vccd1 FuI._028_ sky130_fd_sc_hd__nand2_1
XANTENNA__08951__A _01394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11423_ _04063_ _04062_ _04061_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__a21bo_1
XFILLER_172_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07779__B1 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10378__A2 _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _04121_ _04123_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__a21o_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _02992_ _02993_ _02978_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11285_ _03913_ _03910_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__or4bb_2
XFILLER_3_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ _05853_ _03680_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__or2b_1
X_13024_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__inv_2
XFILLER_140_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3740_ MuI.a_operand\[16\] vssd1 vssd1 vccd1 vccd1 MuI._2840_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12412__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _02808_ _04800_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__and2b_1
XFILLER_20_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3671_ MuI._2583_ MuI._2594_ MuI._2715_ MuI._2726_ vssd1 vssd1 vccd1 vccd1 MuI._2736_
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10098_ _04380_ _02496_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__or2b_1
XFILLER_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5410_ MuI._0100_ MuI._3268_ vssd1 vssd1 vccd1 vccd1 MuI._1194_ sky130_fd_sc_hd__nand2_1
XMuI._6390_ MuI._1966_ MuI._1969_ vssd1 vssd1 vccd1 vccd1 MuI._2272_ sky130_fd_sc_hd__and2_1
XFILLER_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5341_ MuI._1116_ MuI._1117_ vssd1 vssd1 vccd1 vccd1 MuI._1118_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._6046__B MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1215_ AuI._0344_ AuI._0413_ vssd1 vssd1 vccd1 vccd1 AuI._0419_ sky130_fd_sc_hd__and2_1
XFILLER_90_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12648__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5272_ MuI._1039_ MuI._1040_ MuI._1038_ vssd1 vssd1 vccd1 vccd1 MuI._1042_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12808_ _02805_ _05686_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__or2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1146_ AuI._0330_ AuI._0352_ AuI._0231_ AuI._0353_ AuI._0262_ vssd1 vssd1 vccd1
+ vccd1 AuI._0354_ sky130_fd_sc_hd__a311o_1
XFILLER_22_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4223_ MuI._3206_ MuI._3208_ vssd1 vssd1 vccd1 vccd1 MuI._3323_ sky130_fd_sc_hd__nor2_1
XFILLER_188_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12739_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__nand2_1
XAuI._1077_ AuI._0246_ vssd1 vssd1 vccd1 vccd1 AuI._0288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09379__D net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4154_ MuI._3233_ MuI._3253_ vssd1 vssd1 vccd1 vccd1 MuI._3254_ sky130_fd_sc_hd__or2_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4085_ MuI._2880_ vssd1 vssd1 vccd1 vccd1 MuI._3185_ sky130_fd_sc_hd__clkbuf_4
XFILLER_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__B2 _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07477__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5406__A MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5354__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _02609_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__xnor2_2
XFILLER_132_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._747__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08901_ _01349_ _01350_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__nor2_1
XMuI._4987_ MuI._0642_ MuI._0728_ vssd1 vssd1 vccd1 vccd1 MuI._0729_ sky130_fd_sc_hd__nor2_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09881_ _02531_ _02535_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__o21a_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A2 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5106__B1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3938_ MuI._2962_ MuI._2964_ vssd1 vssd1 vccd1 vccd1 MuI._3038_ sky130_fd_sc_hd__nand2_1
XMuI._6726_ MuI._2632_ MuI._2636_ MuI._2641_ vssd1 vssd1 vccd1 vccd1 MuI._2642_ sky130_fd_sc_hd__and3_1
XANTENNA__08734__A2 _01350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08832_ _06548_ _04896_ _04961_ _02291_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22oi_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10541__A2 _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6657_ MuI._2542_ MuI._2565_ MuI._2513_ vssd1 vssd1 vccd1 vccd1 MuI._2566_ sky130_fd_sc_hd__o21a_1
XFILLER_100_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3869_ MuI._2964_ MuI._2965_ MuI._2968_ vssd1 vssd1 vccd1 vccd1 MuI._2969_ sky130_fd_sc_hd__a21o_1
XFILLER_211_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08763_ _01372_ _01379_ _01380_ _01365_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__o211ai_4
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12818__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6237__A MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5779__C MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12818__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5608_ MuI._1397_ MuI._1411_ vssd1 vssd1 vccd1 vccd1 MuI._1412_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._5141__A MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6588_ MuI.a_operand\[23\] MuI._2487_ MuI._0317_ MuI._0295_ vssd1 vssd1 vccd1
+ vccd1 MuI._2490_ sky130_fd_sc_hd__o211a_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07714_ _00328_ _00329_ _00330_ _00331_ vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__a211oi_2
XFILLER_72_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08694_ _01310_ _01309_ _01308_ _01304_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o211a_1
XFILLER_66_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5539_ MuI._3185_ MuI._0110_ MuI.a_operand\[1\] MuI._2892_ vssd1 vssd1 vccd1
+ vccd1 MuI._1336_ sky130_fd_sc_hd__a22o_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07645_ _00262_ _04369_ _00080_ _00087_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__o2bb2a_1
XAuI.pe._419_ AuI.pe.significand\[19\] vssd1 vssd1 vccd1 vccd1 AuI.pe._386_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07576_ _06681_ _00001_ _00003_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__a21bo_1
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09447__B1 _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _02096_ net116 net8 _04767_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__and4_1
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3840__B1 MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0849__B2 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _01855_ _01856_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__o22ai_2
XFILLER_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4396__A1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4396__B2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _01775_ _01782_ _01783_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__and3_1
XANTENNA__09586__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10806__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _00430_ _00433_ _00744_ _00745_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a211o_1
XFILLER_181_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1435__B AuI._0506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _00676_ _04176_ _04240_ _00506_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22oi_1
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11070_ _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__and2b_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1026__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 ALU_Output[19] sky130_fd_sc_hd__buf_2
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10021_ _02676_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nor2_1
XANTENNA__08725__A2 _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__C _01266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ _04786_ _04787_ _04788_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__or3_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10296__A1 _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10923_ _03657_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nand2_1
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1000_ AuI._0157_ AuI._0211_ vssd1 vssd1 vccd1 vccd1 AuI._0212_ sky130_fd_sc_hd__nand2_2
XANTENNA__08665__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10854_ _03582_ _03583_ _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and3_1
XFILLER_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3831__B1 MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _03831_ _04197_ _03353_ _03351_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a31o_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12524_ _05382_ _02900_ _04635_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ _05168_ _05169_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__and2_1
X_11406_ _06428_ _04156_ _04173_ _04180_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__o211ai_4
XANTENNA__07297__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08413__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__B1 _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12386_ _05090_ _05091_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08413__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4910_ MuI._0639_ MuI._0643_ vssd1 vssd1 vccd1 vccd1 MuI._0644_ sky130_fd_sc_hd__xnor2_2
XFILLER_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5890_ MuI._1653_ MuI._1658_ vssd1 vssd1 vccd1 vccd1 MuI._1722_ sky130_fd_sc_hd__nand2_1
XFILLER_141_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ _06429_ _04531_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__and2_2
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._770_ AuI.pe._295_ AuI.pe._313_ vssd1 vssd1 vccd1 vccd1 AuI.pe._314_ sky130_fd_sc_hd__or2_1
XFILLER_107_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4841_ MuI._0566_ MuI._0567_ vssd1 vssd1 vccd1 vccd1 MuI._0568_ sky130_fd_sc_hd__nor2_1
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output77_A net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1017__A1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ _04029_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__nor2_1
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4772_ MuI._0301_ MuI._0302_ MuI._0324_ vssd1 vssd1 vccd1 vccd1 MuI._0492_ sky130_fd_sc_hd__o21a_1
X_13007_ _05803_ _05819_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__or2b_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08716__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ _03067_ _05134_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__and2b_1
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11199_ _03955_ _03953_ _03954_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__nand3_1
XMuI._6511_ MuI._2401_ MuI._2402_ MuI._2404_ vssd1 vssd1 vccd1 vccd1 MuI._2405_ sky130_fd_sc_hd__o21a_1
XMuI._3723_ MuI._2820_ MuI._2822_ vssd1 vssd1 vccd1 vccd1 MuI._2823_ sky130_fd_sc_hd__nor2_1
XFILLER_121_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6442_ MuI._2283_ MuI._2294_ MuI._2293_ vssd1 vssd1 vccd1 vccd1 MuI._2329_ sky130_fd_sc_hd__o21a_1
XFILLER_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3654_ MuI._1296_ vssd1 vssd1 vccd1 vccd1 MuI._2550_ sky130_fd_sc_hd__buf_2
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08856__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6373_ MuI._0867_ MuI._2682_ MuI._2087_ MuI._2089_ vssd1 vssd1 vccd1 vccd1 MuI._2254_
+ sky130_fd_sc_hd__o2bb2a_1
XMuI._3585_ MuI.b_operand\[15\] vssd1 vssd1 vccd1 vccd1 MuI._1791_ sky130_fd_sc_hd__buf_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5324_ MuI._1090_ MuI._1097_ MuI._1099_ vssd1 vssd1 vccd1 vccd1 MuI._1100_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07430_ _00030_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__buf_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12097__B _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5255_ MuI._1017_ MuI._1022_ MuI._1023_ vssd1 vssd1 vccd1 vccd1 MuI._1024_ sky130_fd_sc_hd__nand3_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07361_ _02377_ _06546_ _06550_ _06549_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a31o_1
XAuI._1129_ AuI._0223_ AuI._0199_ AuI._0200_ AuI._0284_ AuI._0208_ vssd1 vssd1 vccd1
+ vccd1 AuI._0338_ sky130_fd_sc_hd__a41o_1
XMuI._4206_ MuI.b_operand\[4\] vssd1 vssd1 vccd1 vccd1 MuI._3306_ sky130_fd_sc_hd__clkbuf_4
X_09100_ _01714_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or2b_1
XFILLER_31_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5186_ MuI._0930_ MuI._0931_ MuI._0946_ vssd1 vssd1 vccd1 vccd1 MuI._0948_ sky130_fd_sc_hd__nand3_1
X_07292_ net122 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__buf_4
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4137_ MuI._0735_ MuI._2813_ MuI._2352_ MuI._2374_ vssd1 vssd1 vccd1 vccd1 MuI._3237_
+ sky130_fd_sc_hd__and4_1
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ _01256_ _01257_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07919__B _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10626__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4068_ MuI._3165_ MuI._3167_ vssd1 vssd1 vccd1 vccd1 MuI._3168_ sky130_fd_sc_hd__xor2_2
XFILLER_129_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__D _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07000__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12841__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4397__D MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ _02592_ _02594_ _02037_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a21oi_1
XANTENNA_AuI._1008__A1 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11457__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09864_ _02488_ _02489_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a21oi_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6709_ MuI._2366_ MuI._2618_ vssd1 vssd1 vccd1 vccd1 MuI._2623_ sky130_fd_sc_hd__or2b_1
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08815_ _03110_ _03906_ _03993_ _03067_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__a22o_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _02322_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__xnor2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _01358_ _01363_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13464__A1 _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__B2 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08766__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07670__A _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6117__D MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _01291_ _01292_ _01294_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__nand3_1
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08485__B _01102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07628_ _00235_ _00245_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__xnor2_2
XFILLER_54_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07559_ _02420_ _06513_ _05434_ _06466_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__nand4_1
XFILLER_195_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ _03180_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__xnor2_2
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07446__A2 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09840__B1 _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09229_ _01676_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__xor2_2
XFILLER_127_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__B _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06733__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _06442_ _00423_ _00002_ _03550_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a22oi_2
XFILLER_135_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3592__A2 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5046__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _02848_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__nand2_1
XFILLER_123_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11950__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ _03871_ _03872_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__xnor2_4
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4100__D MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11053_ _03796_ _03797_ _03779_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a21o_1
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1480_ AuI._0636_ AuI._0665_ vssd1 vssd1 vccd1 vccd1 AuI._0666_ sky130_fd_sc_hd__or2_1
XFILLER_150_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10004_ _01868_ _01872_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__nand2_1
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5097__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08098__D _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12258__A2 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07580__A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _06610_ _05831_ _04656_ _04655_ _05959_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__a32o_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _03594_ _03595_ _03639_ _03640_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__o22a_1
XANTENNA_MuI._3948__B MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__D net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A1 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13207__A1 _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _04694_ _04695_ _04510_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__B2 _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ _03383_ _03385_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__nand2_1
XFILLER_198_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5040_ MuI._0148_ MuI._0281_ vssd1 vssd1 vccd1 vccd1 MuI._0787_ sky130_fd_sc_hd__nor2_1
XFILLER_9_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06924__A _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _02351_ _02745_ _02945_ _04068_ _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a221o_1
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12507_ MuI.result\[16\] _02738_ _04011_ _05363_ _05364_ vssd1 vssd1 vccd1 vccd1
+ _05365_ sky130_fd_sc_hd__a221o_1
XFILLER_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _02750_ _02814_ _06390_ _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__a31o_1
X_10699_ net121 _03047_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__nand2_1
XANTENNA__12718__B1 _05577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _05208_ _05207_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__or2b_1
XANTENNA__07458__C net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12194__A1 _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5942_ MuI._1773_ MuI._1774_ MuI._1777_ MuI._1778_ vssd1 vssd1 vccd1 vccd1 MuI._1779_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12083__D _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12369_ _03798_ _04983_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__nand2_1
XFILLER_181_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._822_ AuI.operand_a\[27\] AuI.pe._197_ vssd1 vssd1 vccd1 vccd1 AuI.pe._360_
+ sky130_fd_sc_hd__xnor2_2
XMuI._5873_ MuI._1700_ MuI._1701_ MuI._1627_ MuI._1629_ vssd1 vssd1 vccd1 vccd1 MuI._1704_
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4824_ MuI._0419_ MuI._0546_ vssd1 vssd1 vccd1 vccd1 MuI._0550_ sky130_fd_sc_hd__xor2_1
XAuI.pe._753_ AuI.pe.significand\[2\] AuI.pe.significand\[3\] AuI.pe._013_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._297_ sky130_fd_sc_hd__or3b_1
X_06930_ _04671_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__and3_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10181__A _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4755_ MuI._0336_ MuI._0338_ vssd1 vssd1 vccd1 vccd1 MuI._0474_ sky130_fd_sc_hd__or2_1
XAuI.pe._684_ AuI.pe._158_ AuI.pe._002_ AuI.pe._053_ AuI.pe._170_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._232_ sky130_fd_sc_hd__a22o_1
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5403__B MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4945__D MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _03928_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__and3_1
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3706_ MuI._2780_ MuI._2795_ MuI._2805_ vssd1 vssd1 vccd1 vccd1 MuI._2806_ sky130_fd_sc_hd__a21o_1
XANTENNA__11427__D _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _02539_ _06613_ _01217_ _01215_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__a31o_1
XFILLER_209_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4686_ MuI._0396_ MuI._0397_ vssd1 vssd1 vccd1 vccd1 MuI._0398_ sky130_fd_sc_hd__or2b_1
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _02211_ _02212_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nor3_1
X_06792_ _03174_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__and3_1
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0879__B_N net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6425_ MuI._1941_ MuI._1955_ vssd1 vssd1 vccd1 vccd1 MuI._2311_ sky130_fd_sc_hd__or2_1
XMuI._3637_ MuI._2352_ vssd1 vssd1 vccd1 vccd1 MuI._2363_ sky130_fd_sc_hd__buf_2
XFILLER_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08531_ _03335_ _03884_ _01145_ _01148_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__and4_1
XANTENNA__10234__A_N _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__C _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6356_ MuI._2202_ MuI._2191_ MuI._2234_ vssd1 vssd1 vccd1 vccd1 MuI._2235_ sky130_fd_sc_hd__o21a_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3568_ MuI._0757_ MuI._0889_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._1604_ sky130_fd_sc_hd__nand3b_1
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08736__D _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _00046_ _00074_ _00090_ _00049_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._6588__A2 MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5307_ MuI._1073_ MuI._1079_ MuI._1080_ vssd1 vssd1 vccd1 vccd1 MuI._1081_ sky130_fd_sc_hd__o21a_1
XANTENNA_AuI._0921__A0 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6287_ MuI._2914_ MuI._0460_ MuI._2122_ MuI._2120_ MuI._2849_ vssd1 vssd1 vccd1
+ vccd1 MuI._2159_ sky130_fd_sc_hd__a32o_1
XFILLER_51_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07413_ _00028_ _00029_ _00030_ _04703_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__and4_1
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3499_ MuI._0823_ MuI._0834_ vssd1 vssd1 vccd1 vccd1 MuI._0845_ sky130_fd_sc_hd__or2_1
X_08393_ _00842_ _00841_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4035__A MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5238_ MuI._2918_ MuI._0304_ MuI._0110_ MuI._2799_ vssd1 vssd1 vccd1 vccd1 MuI._1005_
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07344_ _02205_ net129 net128 _06534_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a22oi_2
XFILLER_195_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09848__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3874__A MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5169_ MuI._0926_ MuI._0927_ MuI._0883_ MuI._0895_ vssd1 vssd1 vccd1 vccd1 MuI._0929_
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07275_ _06511_ _06533_ _06574_ _06575_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a211o_2
XFILLER_164_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ _01630_ _01629_ _01628_ _01537_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__o211a_1
XFILLER_164_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11392__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07665__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07600__A2 _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13134__B1 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ _02347_ _02394_ _02443_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__and3_1
XFILLER_104_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12488__A2 _05341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10522__C _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08199__C _00663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09847_ _02345_ _03873_ _03971_ _02302_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07364__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11160__A2 _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11915__A _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _02345_ _02409_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__and2_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5484__C1 MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _01345_ _01346_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__nand2_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11999__A1 _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11740_ _04537_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__and3_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4590__D MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _04446_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__and3_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _06322_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__xnor2_1
X_10622_ _03176_ _03175_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__or2b_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11215__A3 _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11620__B1 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ _06224_ _06251_ _06250_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__a21o_1
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ _03258_ _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__xor2_1
XAuI._0980_ AuI._0190_ AuI._0191_ vssd1 vssd1 vccd1 vccd1 AuI._0192_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._6160__A MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _06179_ _06180_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__nor2_1
X_10484_ _03186_ _03183_ _03184_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__nand3b_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12176__B2 AuI.result\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _00132_ _00163_ _00385_ _00133_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a22o_1
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10726__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1601_ AuI._0693_ AuI._0767_ AuI._0772_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0773_
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12154_ _04984_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nor2_1
XFILLER_123_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _02757_ _03854_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__or2_1
XAuI._1532_ AuI._0708_ AuI._0705_ AuI._0714_ AuI._0715_ vssd1 vssd1 vccd1 vccd1 AuI.result\[2\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12085_ _04908_ _04909_ _00058_ _05767_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__and4bb_1
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3868__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1463_ AuI._0376_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0649_ sky130_fd_sc_hd__or2_1
X_11036_ _02754_ _02797_ _00398_ _03424_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and4_1
XFILLER_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._580__B2 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4540_ MuI._0230_ MuI._0233_ MuI._0235_ vssd1 vssd1 vccd1 vccd1 MuI._0237_ sky130_fd_sc_hd__nor3_1
XFILLER_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1394_ AuI._0576_ AuI._0583_ vssd1 vssd1 vccd1 vccd1 AuI._0584_ sky130_fd_sc_hd__nand2_1
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4471_ MuI._0156_ MuI._0159_ vssd1 vssd1 vccd1 vccd1 MuI._0161_ sky130_fd_sc_hd__and2_1
XFILLER_92_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6210_ MuI._2063_ MuI._2072_ MuI._2071_ vssd1 vssd1 vccd1 vccd1 MuI._2074_ sky130_fd_sc_hd__a21o_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _05793_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__nand2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08304__B1 _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3678__B MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ _04751_ _04752_ _04593_ _04595_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__o211a_1
XFILLER_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6141_ MuI._3157_ MuI._3179_ MuI._1997_ vssd1 vssd1 vccd1 vccd1 MuI._1998_ sky130_fd_sc_hd__o21ba_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11869_ _03271_ _06562_ _00530_ _03217_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a22o_1
XANTENNA__13481__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6072_ MuI._1873_ MuI._1876_ MuI._1874_ vssd1 vssd1 vccd1 vccd1 MuI._1922_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12403__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5023_ MuI._0765_ MuI._0766_ MuI._0737_ MuI._0767_ vssd1 vssd1 vccd1 vccd1 MuI._0769_
+ sky130_fd_sc_hd__and4b_1
XFILLER_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07830__A2 _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11914__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5925_ MuI._1712_ MuI._1760_ vssd1 vssd1 vccd1 vccd1 MuI._1761_ sky130_fd_sc_hd__or2_1
XFILLER_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11719__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._805_ AuI.pe._342_ AuI.pe._343_ AuI.operand_a\[26\] AuI.pe._333_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._344_ sky130_fd_sc_hd__and4bb_1
XFILLER_88_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5856_ MuI._1613_ MuI._1619_ MuI._1612_ vssd1 vssd1 vccd1 vccd1 MuI._1685_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12541__D _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07962_ _00570_ _00577_ _00578_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._736_ AuI.pe._385_ AuI.pe._384_ AuI.pe._022_ vssd1 vssd1 vccd1 vccd1 AuI.pe._281_
+ sky130_fd_sc_hd__a21o_1
XMuI._4807_ MuI._0530_ MuI._0399_ vssd1 vssd1 vccd1 vccd1 MuI._0531_ sky130_fd_sc_hd__xnor2_1
X_09701_ _02341_ _02343_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__or2_1
X_06913_ _04489_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[8\] sky130_fd_sc_hd__dlymetal6s2s_1
XMuI._5787_ MuI._0743_ MuI._0741_ MuI._0742_ vssd1 vssd1 vccd1 vccd1 MuI._1609_ sky130_fd_sc_hd__or3_1
XFILLER_68_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07893_ _00509_ _00510_ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__nor2_1
XAuI.pe._667_ AuI.pe._013_ AuI.pe.significand\[7\] AuI.pe._197_ AuI.pe._150_ AuI.pe._062_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._216_ sky130_fd_sc_hd__a32o_1
XMuI._4738_ MuI._0440_ MuI._0441_ MuI._0454_ vssd1 vssd1 vccd1 vccd1 MuI._0455_ sky130_fd_sc_hd__and3_1
X_09632_ _06503_ _06504_ _00271_ _04229_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__and4_1
XANTENNA__11735__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _03744_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06829__A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4669_ MuI._0376_ MuI._0377_ MuI._1461_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0379_
+ sky130_fd_sc_hd__and4bb_1
XAuI.pe._598_ AuI.pe.significand\[12\] AuI.pe._025_ AuI.pe._036_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._152_ sky130_fd_sc_hd__a21o_1
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09563_ _02099_ _02098_ _02097_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__o21ai_1
XFILLER_71_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06775_ _03002_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__buf_4
XFILLER_82_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6245__A MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6408_ MuI._2093_ MuI._2096_ MuI._2094_ vssd1 vssd1 vccd1 vccd1 MuI._2292_ sky130_fd_sc_hd__o21ba_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _01129_ _01130_ _01125_ _01126_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__o211a_1
XANTENNA_MuI._3588__B MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09494_ _02117_ _02119_ _02105_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a21o_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6339_ MuI._2170_ MuI._2173_ vssd1 vssd1 vccd1 vccd1 MuI._2216_ sky130_fd_sc_hd__nor2_1
XFILLER_196_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _01060_ _01061_ _01056_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__a21o_1
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12566__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ net106 _06604_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__nand2_1
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._080_ FuI.a_operand\[23\] FuI._044_ FuI._039_ net104 vssd1 vssd1 vccd1 vccd1
+ FuI._045_ sky130_fd_sc_hd__and4b_1
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07327_ _06619_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6194__B1 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09875__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ _02377_ _06477_ _06482_ _06481_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__a31o_1
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3547__A2 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07189_ _06488_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nand2_1
XFILLER_145_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10814__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13421__B_N _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3770__C MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__C _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1386__A0 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11133__A2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _05795_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__xor2_1
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06739__A _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12841_ _06429_ _05391_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__nand2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6155__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3498__B MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _05646_ _05647_ _05508_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o21a_1
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _04518_ _04519_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a21o_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _04206_ _04215_ _04214_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a21o_1
XANTENNA__09488__C _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10708__B _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _04122_ _02302_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__and2b_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11585_ _04371_ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__and2_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1310__B1 AuI._0506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ _03755_ _05842_ _06233_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10536_ _03073_ _03075_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand2_1
XFILLER_183_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0963_ AuI._0174_ vssd1 vssd1 vccd1 vccd1 AuI._0175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12923__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13255_ _06130_ _06131_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__nand2_1
X_10467_ _03167_ _03165_ _03166_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__nand3_2
XAuI._0894_ net57 AuI._0112_ AuI._0113_ vssd1 vssd1 vccd1 vccd1 AuI._0114_ sky130_fd_sc_hd__o21ai_1
XMuI._3971_ MuI._3064_ MuI._3070_ vssd1 vssd1 vccd1 vccd1 MuI._3071_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13100__A _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ _00029_ _00153_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and2_1
XANTENNA__09565__A2 _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13186_ _03489_ _06081_ _06082_ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a31o_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _03080_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__xnor2_2
XMuI._5710_ MuI._1522_ MuI._1523_ vssd1 vssd1 vccd1 vccd1 MuI._1524_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6690_ MuI._0793_ MuI._1841_ MuI._2004_ vssd1 vssd1 vccd1 vccd1 MuI._2602_ sky130_fd_sc_hd__a21boi_1
XFILLER_123_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ _04836_ _04838_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nand2_1
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__D _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5641_ MuI._1370_ MuI._1401_ vssd1 vssd1 vccd1 vccd1 MuI._1448_ sky130_fd_sc_hd__nand2_1
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._553__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1515_ AuI._0606_ AuI._0694_ AuI._0696_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[0\]
+ sky130_fd_sc_hd__o211a_1
X_12068_ _04892_ _02893_ _02926_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__mux2_1
XAuI.pe._521_ AuI.pe.significand\[3\] AuI.pe._050_ AuI.pe._042_ AuI.pe._056_ AuI.pe._080_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._081_ sky130_fd_sc_hd__a221o_1
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5572_ MuI._1331_ MuI._1332_ MuI._1371_ MuI._1294_ vssd1 vssd1 vccd1 vccd1 MuI._1372_
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11019_ _00086_ _00081_ _06623_ _06517_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nand4_1
XAuI._1446_ AuI._0473_ AuI._0477_ vssd1 vssd1 vccd1 vccd1 AuI._0632_ sky130_fd_sc_hd__nor2_1
XMuI._4523_ MuI._0216_ MuI._0217_ MuI._1263_ MuI._0101_ vssd1 vssd1 vccd1 vccd1 MuI._0219_
+ sky130_fd_sc_hd__and4bb_1
XAuI.pe._452_ AuI.pe._377_ AuI.pe._381_ AuI.pe._398_ AuI.pe._018_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._019_ sky130_fd_sc_hd__and4_1
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3689__A MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1377_ AuI._0567_ AuI._0568_ vssd1 vssd1 vccd1 vccd1 AuI._0569_ sky130_fd_sc_hd__or2_2
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4454_ MuI._0132_ MuI._0133_ MuI._0142_ vssd1 vssd1 vccd1 vccd1 MuI._0143_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4385_ MuI._3336_ MuI._0067_ vssd1 vssd1 vccd1 vccd1 MuI._0068_ sky130_fd_sc_hd__or2_1
XMuI._6124_ MuI._1977_ MuI._1979_ vssd1 vssd1 vccd1 vccd1 MuI._1980_ sky130_fd_sc_hd__nor2_1
XFILLER_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._608__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08230_ _00635_ _00636_ _00637_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__and3_1
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6055_ MuI._1883_ MuI._1903_ vssd1 vssd1 vccd1 vccd1 MuI._1904_ sky130_fd_sc_hd__xor2_1
XANTENNA__12388__A1 _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3777__A2 MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08161_ _00776_ _00777_ _00772_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__a21o_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5006_ MuI._0747_ MuI._0748_ MuI._0749_ vssd1 vssd1 vccd1 vccd1 MuI._0750_ sky130_fd_sc_hd__nand3_2
X_07112_ _05595_ _06414_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08092_ _00691_ _00709_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4726__A1 MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _05884_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__buf_4
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10634__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout109_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._792__A1 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5908_ MuI._1675_ MuI._1677_ vssd1 vssd1 vccd1 vccd1 MuI._1742_ sky130_fd_sc_hd__and2_1
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08994_ _01372_ _01379_ _01380_ _01365_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__o211a_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5839_ MuI._1565_ MuI._1469_ MuI._1468_ MuI._1467_ vssd1 vssd1 vccd1 vccd1 MuI._1666_
+ sky130_fd_sc_hd__and4b_1
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07945_ _00070_ _00071_ _00105_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__nor3_2
XAuI.pe._719_ AuI.pe._158_ AuI.pe._399_ AuI.pe._053_ AuI.pe._201_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._265_ sky130_fd_sc_hd__a22o_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11115__A2 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07662__B _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07876_ _00491_ _00492_ _00485_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a21o_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09615_ _02242_ _02250_ _02251_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a21bo_1
X_06827_ _03561_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__and3_1
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09546_ _06513_ _04100_ _04165_ _02420_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
X_06758_ _02819_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[13\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__08774__A _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11823__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _06545_ _00259_ _02043_ _02044_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__o2bb2a_1
X_06689_ _02053_ _02075_ vssd1 vssd1 vccd1 vccd1 AuI.AddBar_Sub sky130_fd_sc_hd__nand2_2
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ _01043_ _01044_ _01045_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__nand3_1
XFILLER_180_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1438__B AuI._0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._132_ FuI._016_ net138 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[3\] sky130_fd_sc_hd__dlxtn_1
XFILLER_200_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08047__A2 _00663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _00971_ _00972_ _00976_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__a21o_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11370_ _03989_ _03991_ _04140_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__a211oi_4
XFILLER_192_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10321_ _03013_ _04983_ _03009_ _03010_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nand4_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _05923_ _05924_ _05925_ _05926_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a221o_1
X_10252_ _02730_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__A1 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__B2 _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _04994_ _02970_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__and2b_1
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1071__A2 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5142__A1 MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5142__B2 MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._535__B2 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A b_operand[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1300_ AuI._0487_ vssd1 vssd1 vccd1 vccd1 AuI._0498_ sky130_fd_sc_hd__buf_2
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1231_ AuI._0433_ AuI._0434_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[8\]
+ sky130_fd_sc_hd__nor2_2
XANTENNA__07291__C _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12824_ _05701_ _05703_ _05697_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__o21ai_1
XAuI._1162_ AuI._0274_ AuI._0268_ AuI._0368_ AuI._0276_ vssd1 vssd1 vccd1 vccd1 AuI._0369_
+ sky130_fd_sc_hd__a211o_1
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1093_ AuI._0302_ AuI._0303_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[1\]
+ sky130_fd_sc_hd__nor2_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _00676_ _05445_ _05509_ _00506_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a22oi_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4170_ MuI._3263_ MuI._3267_ MuI._3269_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._3270_
+ sky130_fd_sc_hd__o211a_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11706_ _05895_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3956__B MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4405__B1 MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _05492_ _05466_ _05555_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o211ai_4
XANTENNA_AuI._0885__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4956__A1 MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5229__A MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4956__B2 MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11637_ _04269_ _04287_ _04288_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._3675__C MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11568_ FuI.Integer\[9\] _06045_ _02718_ _04607_ vssd1 vssd1 vccd1 vccd1 _04354_
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06932__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4708__A1 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3972__A MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4708__B2 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13307_ _02751_ _06162_ _06163_ _06217_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__a31o_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10519_ _03223_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nor2_1
XFILLER_183_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0946_ net56 net131 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0158_ sky130_fd_sc_hd__mux2_1
X_11499_ _04278_ _04279_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a21o_1
XMuI._6811_ MuI._2734_ vssd1 vssd1 vccd1 vccd1 MuI._2735_ sky130_fd_sc_hd__buf_2
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ FuI.Integer\[25\] _06045_ _02744_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11269__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0877_ net55 net23 vssd1 vssd1 vccd1 vccd1 AuI._0097_ sky130_fd_sc_hd__xor2_2
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6742_ MuI._2475_ MuI._2658_ vssd1 vssd1 vccd1 vccd1 MuI._2659_ sky130_fd_sc_hd__nor2_1
XMuI._3954_ MuI._3046_ MuI._3047_ MuI._3052_ vssd1 vssd1 vccd1 vccd1 MuI._3054_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08210__A2 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _04678_ _05052_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__a21o_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5133__A1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3885_ MuI._2840_ MuI._2802_ MuI._2649_ MuI._2843_ vssd1 vssd1 vccd1 vccd1 MuI._2985_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._5133__B2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6673_ MuI._0282_ MuI._2581_ vssd1 vssd1 vccd1 vccd1 MuI._2584_ sky130_fd_sc_hd__nand2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5624_ MuI._1401_ MuI._1409_ MuI._1429_ vssd1 vssd1 vccd1 vccd1 MuI._1430_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11285__A _03913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07730_ _00345_ _04186_ _00346_ _00347_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__nand4_1
XFILLER_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._504_ AuI.pe.significand\[5\] AuI.pe.significand\[4\] AuI.pe._049_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._065_ sky130_fd_sc_hd__or3_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5555_ MuI._1350_ MuI._1352_ MuI._1353_ vssd1 vssd1 vccd1 vccd1 MuI._1354_ sky130_fd_sc_hd__o21bai_1
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1429_ AuI._0557_ AuI._0560_ vssd1 vssd1 vccd1 vccd1 AuI._0615_ sky130_fd_sc_hd__or2b_1
X_07661_ net54 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._435_ AuI.pe._001_ vssd1 vssd1 vccd1 vccd1 AuI.pe._002_ sky130_fd_sc_hd__buf_2
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4506_ MuI._0176_ MuI._0197_ MuI._0199_ vssd1 vssd1 vccd1 vccd1 MuI._0200_ sky130_fd_sc_hd__a21oi_1
X_09400_ _01946_ _01949_ _01948_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__o21ai_2
XFILLER_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5486_ MuI._1276_ MuI._1277_ vssd1 vssd1 vccd1 vccd1 MuI._1278_ sky130_fd_sc_hd__or2_1
XANTENNA__12058__B1 _01233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4644__B1 MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ _00186_ _00187_ _00209_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__o21ai_2
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4437_ MuI._3378_ MuI._0122_ MuI._0121_ MuI._0071_ vssd1 vssd1 vccd1 vccd1 MuI._0124_
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ _01945_ _01944_ _01943_ _01939_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o211a_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4368_ MuI._0037_ MuI._0047_ MuI._0048_ vssd1 vssd1 vccd1 vccd1 MuI._0049_ sky130_fd_sc_hd__a21oi_2
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _01878_ _01879_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__and2_1
XFILLER_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6107_ MuI._1959_ MuI._1878_ MuI._1960_ vssd1 vssd1 vccd1 vccd1 MuI._1961_ sky130_fd_sc_hd__o21bai_1
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6242__B MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08213_ _00825_ _00826_ _00830_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__a21o_1
XANTENNA__07003__A _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4299_ MuI._3263_ MuI._3398_ vssd1 vssd1 vccd1 vccd1 MuI._3399_ sky130_fd_sc_hd__xor2_1
X_09193_ _01755_ _01756_ _01757_ _01735_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6038_ MuI._1884_ vssd1 vssd1 vccd1 vccd1 MuI._1885_ sky130_fd_sc_hd__inv_2
X_08144_ _00759_ _00760_ _00761_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__nand3_2
XANTENNA__07237__B1 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06842__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _00270_ _00093_ _00457_ _00230_ _00036_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a32o_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07026_ _05702_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__buf_2
XFILLER_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._765__B2 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__B _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08737__B1 _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11907__B _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _06491_ _06604_ _06580_ _06492_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a22oi_2
XFILLER_130_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5675__A2 MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07392__B _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07928_ _00414_ _06579_ _04896_ _06580_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__and4_1
XFILLER_69_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07859_ _00441_ _00476_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _03600_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__nor2_1
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08981__A1_N _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _02147_ _02148_ _02157_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__and4bb_1
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11642__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10539__A net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12540_ _03282_ _05702_ _05767_ _03228_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__a22oi_1
XFILLER_185_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08009__A _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0867__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ _05308_ _05324_ _05325_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and3_1
XFILLER_138_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFuI._115_ net105 FuI.a_operand\[29\] FuI.a_operand\[28\] FuI.a_operand\[27\] vssd1
+ vssd1 vccd1 vccd1 FuI._027_ sky130_fd_sc_hd__and4b_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11422_ _04195_ _04193_ _04194_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__nand3_1
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06752__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07779__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07779__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _03885_ _03887_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _02978_ _02992_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__and3_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11284_ _04045_ _04047_ _04028_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__a21o_1
XANTENNA__07286__C _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13023_ _05748_ _05835_ _05837_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__nand3_1
X_10235_ _02917_ _05917_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__or2_1
XFILLER_133_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._508__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10166_ _04800_ _02808_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__or2b_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3670_ MuI._2704_ MuI._2616_ MuI._2649_ MuI._2671_ vssd1 vssd1 vccd1 vccd1 MuI._2726_
+ sky130_fd_sc_hd__and4_1
XFILLER_94_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10097_ _02496_ _04391_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__or2b_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5340_ MuI._1114_ MuI._1115_ MuI._1108_ MuI._1113_ vssd1 vssd1 vccd1 vccd1 MuI._1117_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1214_ AuI._0404_ AuI._0418_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[7\]
+ sky130_fd_sc_hd__xnor2_4
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06927__A _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5271_ MuI._1038_ MuI._1039_ MuI._1040_ vssd1 vssd1 vccd1 vccd1 MuI._1041_ sky130_fd_sc_hd__or3_1
XANTENNA__12648__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3967__A MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _02805_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__nand2_1
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1145_ AuI._0236_ AuI._0241_ AuI._0209_ vssd1 vssd1 vccd1 vccd1 AuI._0353_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4222_ MuI._3319_ MuI._3321_ vssd1 vssd1 vccd1 vccd1 MuI._3322_ sky130_fd_sc_hd__or2b_1
X_10999_ _03588_ _03571_ _03573_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand3_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._692__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05500_ _05506_ _05499_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__a21o_1
XAuI._1076_ AuI._0276_ AuI._0281_ AuI._0286_ AuI._0153_ vssd1 vssd1 vccd1 vccd1 AuI._0287_
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4153_ MuI._3233_ MuI._3234_ MuI._3252_ vssd1 vssd1 vccd1 vccd1 MuI._3253_ sky130_fd_sc_hd__nor3_1
XFILLER_31_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12669_ _05537_ _05535_ _05536_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__nand3_1
XMuI._4084_ MuI._0570_ MuI._2886_ MuI._2882_ MuI._0328_ vssd1 vssd1 vccd1 vccd1 MuI._3184_
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11566__A2 _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5354__A1 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5354__B2 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5406__B MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0929_ AuI._0128_ AuI._0129_ net52 vssd1 vssd1 vccd1 vccd1 AuI._0141_ sky130_fd_sc_hd__a21o_1
XFILLER_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08900_ _01516_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__nor2_1
XFILLER_125_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4986_ MuI._2817_ MuI._0320_ MuI._0640_ MuI._0641_ vssd1 vssd1 vccd1 vccd1 MuI._0728_
+ sky130_fd_sc_hd__o2bb2a_1
X_09880_ _02495_ _02536_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__nor2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5106__A1 MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6725_ MuI._2635_ MuI._2640_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2641_ sky130_fd_sc_hd__mux2_1
XFILLER_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5106__B2 MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3937_ MuI._3035_ MuI._3036_ vssd1 vssd1 vccd1 vccd1 MuI._3037_ sky130_fd_sc_hd__xnor2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _06544_ _06603_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__nand2_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5422__A MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6656_ MuI._2557_ MuI._2564_ MuI._2544_ MuI._2551_ vssd1 vssd1 vccd1 vccd1 MuI._2565_
+ sky130_fd_sc_hd__a211o_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3868_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._2893_ MuI._2967_ vssd1
+ vssd1 vccd1 vccd1 MuI._2968_ sky130_fd_sc_hd__o311a_1
X_08762_ _01342_ _01347_ _01364_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__nand3_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12818__A2 _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5607_ MuI._1393_ MuI._1394_ MuI._1396_ vssd1 vssd1 vccd1 vccd1 MuI._1411_ sky130_fd_sc_hd__o21ba_1
XANTENNA_MuI._6237__B MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5779__D MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07713_ _00286_ _00295_ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__and2b_1
XMuI._3799_ MuI._1032_ MuI._2898_ vssd1 vssd1 vccd1 vccd1 MuI._2899_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5141__B MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6587_ MuI.a_operand\[23\] MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2489_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08693_ _01304_ _01308_ _01309_ _01310_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10610__A_N _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5538_ MuI._2886_ MuI._2882_ MuI._0111_ MuI._0315_ vssd1 vssd1 vccd1 vccd1 MuI._1335_
+ sky130_fd_sc_hd__and4_1
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _00088_ vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__buf_4
XAuI.pe._418_ AuI.pe.significand\[18\] vssd1 vssd1 vccd1 vccd1 AuI.pe._385_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06837__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5469_ MuI._1249_ MuI._1257_ MuI._1258_ vssd1 vssd1 vccd1 vccd1 MuI._1259_ sky130_fd_sc_hd__a21bo_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09447__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _00190_ _00191_ _00189_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09447__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09314_ _00150_ _00032_ _04767_ _06469_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a22oi_2
XFILLER_179_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3840__A1 MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3840__B2 MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0849__A2 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _01860_ _01861_ _01650_ _01857_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__o211a_1
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4396__A2 MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _01789_ _01790_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nand3_1
XANTENNA__13389__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09586__C _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10806__B _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _00725_ _00726_ _00743_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__nor3b_1
XFILLER_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07630__B1 _00246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _03593_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__buf_2
XFILLER_190_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__A1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12506__B2 _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _05520_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 ALU_Output[0] sky130_fd_sc_hd__buf_2
XANTENNA__10517__B1 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10020_ _02662_ _02675_ _02674_ _02671_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a211oi_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11971_ net114 _03047_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__nand2_1
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ _03509_ _03510_ _03656_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nand3_1
XANTENNA__10296__A2 _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06747__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12690__B1 _05559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08665__C _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4084__A1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _03403_ _03401_ _03402_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._4084__B2 MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10269__A _00707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._674__B1 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10784_ _03332_ _03483_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nand2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12523_ _02865_ _05261_ _02864_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a21o_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12454_ _05306_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and2_1
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _02773_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5507__A MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _05087_ _05089_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
XANTENNA__08413__A2 _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__xor2_4
XFILLER_181_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4840_ MuI._0562_ MuI._0565_ vssd1 vssd1 vccd1 vccd1 MuI._0567_ sky130_fd_sc_hd__and2_1
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11267_ _00012_ _00011_ _03425_ _05702_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__and4_1
XFILLER_106_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _05881_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__xnor2_1
XMuI._4771_ MuI._0485_ MuI._0489_ MuI._0490_ MuI._0476_ vssd1 vssd1 vccd1 vccd1 MuI._0491_
+ sky130_fd_sc_hd__o211ai_2
X_10218_ _02849_ _02900_ _02850_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21o_1
XFILLER_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11198_ _03953_ _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__a21o_1
XMuI._6510_ MuI._2121_ MuI._2403_ vssd1 vssd1 vccd1 vccd1 MuI._2404_ sky130_fd_sc_hd__nor2_1
XMuI._3722_ MuI._2820_ MuI._2821_ MuI._0867_ MuI._2385_ vssd1 vssd1 vccd1 vccd1 MuI._2822_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA_MuI._4784__C MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _03561_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__inv_2
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4847__B1 MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3653_ MuI._2451_ vssd1 vssd1 vccd1 vccd1 MuI._2539_ sky130_fd_sc_hd__buf_2
XMuI._6441_ MuI._2320_ MuI._2326_ MuI._2327_ vssd1 vssd1 vccd1 vccd1 MuI._2328_ sky130_fd_sc_hd__nand3_1
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08856__B _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6372_ MuI._2245_ MuI._2246_ MuI._2249_ vssd1 vssd1 vccd1 vccd1 MuI._2252_ sky130_fd_sc_hd__and3_1
XMuI._3584_ MuI._1538_ MuI._1769_ vssd1 vssd1 vccd1 vccd1 MuI._1780_ sky130_fd_sc_hd__nand2_1
XFILLER_208_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5323_ MuI._1091_ MuI._1092_ MuI._1096_ vssd1 vssd1 vccd1 vccd1 MuI._1099_ sky130_fd_sc_hd__nand3_1
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1089__A AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10179__A _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5254_ MuI._1019_ MuI._1020_ MuI._1018_ vssd1 vssd1 vccd1 vccd1 MuI._1023_ sky130_fd_sc_hd__a21bo_1
XFILLER_204_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09968__A _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _06566_ _06567_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nand2_1
XAuI._1128_ AuI._0307_ AuI._0192_ AuI._0277_ vssd1 vssd1 vccd1 vccd1 AuI._0337_ sky130_fd_sc_hd__and3_1
XFILLER_210_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4205_ MuI._3300_ MuI._3298_ vssd1 vssd1 vccd1 vccd1 MuI._3305_ sky130_fd_sc_hd__xor2_2
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5185_ MuI._0930_ MuI._0931_ MuI._0946_ vssd1 vssd1 vccd1 vccd1 MuI._0947_ sky130_fd_sc_hd__a21o_1
XANTENNA__12984__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07291_ _06589_ _06590_ _02712_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__and4bb_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1059_ AuI._0164_ AuI._0169_ AuI._0220_ vssd1 vssd1 vccd1 vccd1 AuI._0270_ sky130_fd_sc_hd__and3_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4136_ MuI._2822_ MuI._3235_ vssd1 vssd1 vccd1 vccd1 MuI._3236_ sky130_fd_sc_hd__nor2_1
X_09030_ _01570_ _01574_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__nand2_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07919__C _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10626__B _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4067_ MuI._3075_ MuI._3166_ vssd1 vssd1 vccd1 vccd1 MuI._3167_ sky130_fd_sc_hd__or2_1
XFILLER_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4321__A MuI._3418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12841__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _02035_ _02036_ _02032_ _02034_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a211o_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4969_ MuI._0693_ MuI._0707_ MuI._0708_ MuI._0646_ vssd1 vssd1 vccd1 vccd1 MuI._0709_
+ sky130_fd_sc_hd__a211o_2
X_09863_ _02450_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__nand2_1
XANTENNA__11457__B _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08112__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6708_ MuI._2619_ vssd1 vssd1 vccd1 vccd1 MuI._2622_ sky130_fd_sc_hd__clkinv_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5152__A MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08814_ _01430_ _01423_ _01429_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nand3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _02347_ _02394_ _02317_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6639_ MuI._1454_ MuI._1456_ vssd1 vssd1 vccd1 vccd1 MuI._2546_ sky130_fd_sc_hd__xnor2_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08745_ _01361_ _01362_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4991__A MuI._0725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13464__A2 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__B net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__B _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08676_ _01218_ _01293_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__xor2_1
XFILLER_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__B _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07627_ _00243_ _00244_ vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__or2b_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5263__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09878__A _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _06513_ _05434_ _06466_ _02420_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__a22o_1
XANTENNA__12424__B1 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09840__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _00057_ _00066_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__or2b_1
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ _01767_ _01844_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a21boi_1
XANTENNA_AuI._1446__B AuI._0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__C _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09159_ net106 _00089_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__nand2_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5046__B MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _02843_ _04883_ _00566_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__o21bai_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ _03722_ _04456_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__and2_2
XFILLER_162_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _03779_ _03796_ _03797_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__nand3_2
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10003_ _01866_ _02667_ _02668_ _02670_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__o211a_1
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input21_A a_operand[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0806__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07580__B _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ _04661_ _04659_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2b_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__A2 _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _03594_ _03595_ _03639_ _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__nor4_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ _04510_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__and3_1
XANTENNA__13207__A2 _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A2 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _03563_ _03564_ _03559_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a21o_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12966__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _02302_ _04133_ _02721_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__o21a_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6203__C1 MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10977__B1 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10727__A _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _02970_ _04994_ _02743_ _02944_ _04929_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__a32o_1
XFILLER_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10186__A_N _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _02741_ _06394_ _06395_ _06396_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a311o_1
X_10698_ _03244_ _03253_ _03252_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__a21bo_1
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10446__B _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07101__A _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5237__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ _05287_ _05288_ _05267_ _05174_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__a211o_1
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07458__D _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5941_ MuI._0733_ MuI._1776_ MuI._1749_ MuI._1775_ vssd1 vssd1 vccd1 vccd1 MuI._1778_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _05213_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._821_ AuI.pe._358_ AuI.pe._359_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[3\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__06940__A _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5872_ MuI._1627_ MuI._1629_ MuI._1700_ MuI._1701_ vssd1 vssd1 vccd1 vccd1 MuI._1702_
+ sky130_fd_sc_hd__o211ai_1
X_11319_ _04085_ _04067_ _04069_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__and3_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10462__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ _05140_ _02898_ _04635_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__mux2_1
XAuI.pe._752_ AuI.pe._013_ AuI.pe._274_ AuI.pe._256_ AuI.pe.significand\[2\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._296_ sky130_fd_sc_hd__a22o_1
XMuI._4823_ MuI._0285_ MuI._0417_ vssd1 vssd1 vccd1 vccd1 MuI._0549_ sky130_fd_sc_hd__xor2_1
XFILLER_141_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09898__A1 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._683_ AuI.pe._145_ AuI.pe._079_ AuI.pe._119_ AuI.pe._102_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._231_ sky130_fd_sc_hd__a22o_1
XFILLER_110_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4754_ MuI._0469_ MuI._0472_ vssd1 vssd1 vccd1 vccd1 MuI._0473_ sky130_fd_sc_hd__or2b_1
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06860_ _03917_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__buf_4
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3705_ MuI._2798_ MuI._2801_ MuI._2804_ vssd1 vssd1 vccd1 vccd1 MuI._2805_ sky130_fd_sc_hd__o21bai_1
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4685_ MuI._0167_ MuI._0179_ vssd1 vssd1 vccd1 vccd1 MuI._0397_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06791_ _02151_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__clkbuf_2
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6424_ MuI._2278_ MuI._2279_ MuI._2281_ vssd1 vssd1 vccd1 vccd1 MuI._2310_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08586__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3636_ MuI._2341_ vssd1 vssd1 vccd1 vccd1 MuI._2352_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ _01146_ _06437_ _06443_ _01147_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__a22o_1
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07921__D _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6355_ MuI._2232_ MuI._2233_ vssd1 vssd1 vccd1 vccd1 MuI._2234_ sky130_fd_sc_hd__nor2_1
XMuI._3567_ MuI._1076_ MuI._1582_ vssd1 vssd1 vccd1 vccd1 MuI._1593_ sky130_fd_sc_hd__xnor2_1
X_08461_ _00028_ _00029_ _04294_ _00072_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__and4_1
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5306_ MuI._0838_ MuI._0839_ vssd1 vssd1 vccd1 vccd1 MuI._1080_ sky130_fd_sc_hd__xnor2_1
X_07412_ net7 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0921__A1 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6286_ MuI._2156_ MuI._2157_ vssd1 vssd1 vccd1 vccd1 MuI._2158_ sky130_fd_sc_hd__xnor2_1
XMuI._3498_ MuI._0636_ MuI._0592_ MuI._0394_ vssd1 vssd1 vccd1 vccd1 MuI._0834_ sky130_fd_sc_hd__and3_1
XFILLER_196_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _00965_ _00966_ _00967_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__o21ba_1
XFILLER_51_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4035__B MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5237_ MuI._2693_ MuI._2638_ MuI._0304_ MuI._0444_ vssd1 vssd1 vccd1 vccd1 MuI._1004_
+ sky130_fd_sc_hd__and4_1
XFILLER_177_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07343_ _02248_ net130 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__nand2_1
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09848__D _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5168_ MuI._0883_ MuI._0895_ MuI._0926_ MuI._0927_ vssd1 vssd1 vccd1 vccd1 MuI._0928_
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_MuI._3874__B MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07274_ _06556_ _06557_ _06573_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__and3_1
XFILLER_176_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4119_ MuI._3216_ MuI._3217_ MuI._3218_ vssd1 vssd1 vccd1 vccd1 MuI._3219_ sky130_fd_sc_hd__o21ba_1
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _01537_ _01628_ _01629_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a211oi_4
XMuI._5099_ MuI._0849_ MuI._0850_ MuI._0848_ vssd1 vssd1 vccd1 vccd1 MuI._0852_ sky130_fd_sc_hd__o21ai_1
XFILLER_164_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13034__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06850__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13134__A1 _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13134__B2 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09915_ _02521_ _02573_ _02574_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a21o_1
XFILLER_160_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10522__D _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _02497_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__or2b_1
XFILLER_112_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__A2 _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07681__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _02371_ _02425_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__or2_1
XANTENNA__11915__B _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5484__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__A2 _06345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06989_ _05305_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__buf_4
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5610__A MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _01336_ _01341_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__xnor2_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__B1 _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08659_ _01135_ _01136_ _01173_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__o21ai_1
XANTENNA_MuI._4226__A MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ _04462_ _04463_ _04283_ _04447_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__a211o_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _03139_ _03179_ _03333_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__o21ai_2
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5539__A1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ _06224_ _06250_ _06251_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__and3_1
XFILLER_210_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5539__B2 MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11620__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _05948_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a21bo_1
XFILLER_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11620__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6160__B MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__C _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _06167_ _06116_ _06178_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and3_1
X_10483_ _03183_ _03184_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12762__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12222_ _00921_ _00132_ _05702_ _03247_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nand4_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06760__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1600_ AuI._0625_ AuI._0771_ vssd1 vssd1 vccd1 vccd1 AuI._0772_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12153_ _04981_ _04982_ _04939_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10282__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11104_ _02757_ _03854_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI._0828__A_N net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._1531_ AuI.pe.Significand\[2\] AuI._0695_ AuI.Exception vssd1 vssd1 vccd1 vccd1
+ AuI._0715_ sky130_fd_sc_hd__o21ba_1
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12084_ _00444_ _05767_ _04908_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11035_ _00011_ _05509_ _05574_ _00012_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a22oi_1
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1462_ AuI._0411_ AuI._0415_ vssd1 vssd1 vccd1 vccd1 AuI._0648_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12884__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1393_ AuI._0389_ AuI._0276_ AuI._0390_ AuI._0422_ vssd1 vssd1 vccd1 vccd1 AuI._0583_
+ sky130_fd_sc_hd__and4_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4470_ MuI._0156_ MuI._0159_ vssd1 vssd1 vccd1 vccd1 MuI._0160_ sky130_fd_sc_hd__nor2_1
XFILLER_94_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12986_ _05796_ _05795_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__or2b_1
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__A1 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__B2 _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _04593_ _04595_ _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a211oi_4
XFILLER_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6140_ MuI._3180_ MuI._2960_ vssd1 vssd1 vccd1 vccd1 MuI._1997_ sky130_fd_sc_hd__and2b_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11868_ _00125_ _00530_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__nand2_2
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06935__A _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6071_ MuI._1919_ MuI._1920_ vssd1 vssd1 vccd1 vccd1 MuI._1921_ sky130_fd_sc_hd__xor2_1
XFILLER_159_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10819_ _03545_ _03543_ _03544_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__nand3_1
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ _04475_ _04497_ _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__o211ai_4
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5022_ MuI._0709_ MuI._0736_ MuI._0725_ MuI._0734_ vssd1 vssd1 vccd1 vccd1 MuI._0767_
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13469_ _06428_ _06362_ _06363_ _06366_ _06384_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__o311ai_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07766__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5924_ MuI._1713_ MuI._1759_ vssd1 vssd1 vccd1 vccd1 MuI._1760_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11914__A2 _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._804_ AuI.pe._392_ AuI.pe._096_ AuI.pe._118_ AuI.pe._150_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._343_ sky130_fd_sc_hd__or4_1
XFILLER_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5855_ MuI._1607_ MuI._1622_ MuI._1623_ vssd1 vssd1 vccd1 vccd1 MuI._1684_ sky130_fd_sc_hd__nand3_1
X_07961_ _00570_ _00577_ _00578_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__a21o_1
XFILLER_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._735_ AuI.pe.significand\[21\] AuI.pe._026_ AuI.pe._002_ AuI.pe._201_ AuI.pe._037_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._280_ sky130_fd_sc_hd__a221o_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4806_ MuI._0396_ MuI._0397_ vssd1 vssd1 vccd1 vccd1 MuI._0530_ sky130_fd_sc_hd__xor2_1
X_09700_ _02219_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__nor2_1
XANTENNA__10201__A_N _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06912_ _04467_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__and3_1
XMuI._5786_ MuI._1524_ MuI._1533_ MuI._1532_ vssd1 vssd1 vccd1 vccd1 MuI._1608_ sky130_fd_sc_hd__a21bo_1
XFILLER_96_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._571__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07892_ _06439_ _04046_ _00507_ _00508_ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08597__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._666_ AuI.pe._059_ AuI.pe._164_ AuI.pe._214_ vssd1 vssd1 vccd1 vccd1 AuI.pe._215_
+ sky130_fd_sc_hd__a21o_1
XMuI._4737_ MuI._0450_ MuI._0453_ vssd1 vssd1 vccd1 vccd1 MuI._0454_ sky130_fd_sc_hd__xor2_1
X_09631_ _02267_ _02268_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__or2_1
XFILLER_110_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__B _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06843_ _03733_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4972__C MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._597_ AuI.pe._062_ AuI.pe._086_ AuI.pe._066_ AuI.pe._089_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._151_ sky130_fd_sc_hd__a22o_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4668_ MuI.b_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._0378_ sky130_fd_sc_hd__clkbuf_4
X_09562_ _02099_ _02097_ _02098_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__or3_1
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06774_ net119 vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__buf_4
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6407_ MuI._2289_ MuI._2290_ vssd1 vssd1 vccd1 vccd1 MuI._2291_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._6245__B MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3619_ MuI._1362_ MuI._1406_ MuI._2154_ vssd1 vssd1 vccd1 vccd1 MuI._2165_ sky130_fd_sc_hd__o21a_1
XANTENNA__07006__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ _01125_ _01126_ _01129_ _01130_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a211oi_4
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4599_ MuI._0300_ MuI._0291_ MuI._0299_ vssd1 vssd1 vccd1 vccd1 MuI._0302_ sky130_fd_sc_hd__and3_1
X_09493_ _02105_ _02117_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__nand3_2
XFILLER_24_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6338_ MuI._1956_ MuI._2214_ vssd1 vssd1 vccd1 vccd1 MuI._2215_ sky130_fd_sc_hd__nor2_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08444_ _01056_ _01060_ _01061_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__nand3_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12566__B _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6269_ MuI._2137_ MuI._2138_ vssd1 vssd1 vccd1 vccd1 MuI._2139_ sky130_fd_sc_hd__xor2_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__B1 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08375_ net107 net66 net133 net13 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__and4_1
XFILLER_177_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07326_ _06621_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07806__B1 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10086__B _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09875__B _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07257_ _02550_ _05198_ _06528_ _06527_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a31o_1
XFILLER_192_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13355__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07188_ net20 vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10814__B _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13107__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3770__D MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__D _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1386__A1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _02450_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__nand2_1
XFILLER_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ _05720_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6155__B MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _05508_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__nor3_2
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _04388_ _04390_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__nand2_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3795__A MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11653_ _04121_ _04126_ _04283_ _04284_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a211oi_2
XFILLER_30_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10277__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09488__D _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _02556_ _02562_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__or2_1
XFILLER_211_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _04225_ _04226_ _04370_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__nand3_1
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ _03755_ _05842_ _06233_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and3_1
XFILLER_128_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ _03241_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__nor2_1
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0962_ AuI._0029_ AuI._0030_ vssd1 vssd1 vccd1 vccd1 AuI._0174_ sky130_fd_sc_hd__nor2_1
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13346__A1 _05700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13254_ _02833_ _06161_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__nand2_1
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10466_ _03165_ _03166_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__a21o_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0893_ net58 net128 vssd1 vssd1 vccd1 vccd1 AuI._0113_ sky130_fd_sc_hd__or2b_1
X_12205_ _02905_ _05959_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__nand2_1
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3970_ MuI._3066_ MuI._3069_ vssd1 vssd1 vccd1 vccd1 MuI._3070_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _06084_ _06088_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__or3_1
X_10397_ _03091_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08773__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ _04963_ _04964_ _04959_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a21o_1
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5696__B1 MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5640_ MuI._1430_ MuI._1445_ MuI._1446_ vssd1 vssd1 vccd1 vccd1 MuI._1447_ sky130_fd_sc_hd__a21o_1
XAuI._1514_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0700_ sky130_fd_sc_hd__buf_2
XFILLER_111_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ _02869_ _04634_ _02870_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__o21bai_1
XAuI.pe._520_ AuI.pe._071_ AuI.pe._026_ AuI.pe._022_ AuI.pe._062_ AuI.pe._037_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._080_ sky130_fd_sc_hd__a221o_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5571_ MuI._1334_ MuI._1370_ vssd1 vssd1 vccd1 vccd1 MuI._1371_ sky130_fd_sc_hd__nor2_1
X_11018_ _00096_ _05101_ _06517_ _00095_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__a22o_1
XAuI._1445_ AuI._0625_ AuI._0626_ vssd1 vssd1 vccd1 vccd1 AuI._0631_ sky130_fd_sc_hd__nand2_1
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._451_ AuI.pe._007_ AuI.pe._012_ AuI.pe._016_ AuI.pe._017_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._018_ sky130_fd_sc_hd__and4bb_1
XFILLER_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4522_ MuI._1802_ MuI._2374_ MuI._3363_ MuI._1307_ vssd1 vssd1 vccd1 vccd1 MuI._0217_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5250__A MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1376_ AuI._0257_ AuI._0565_ AuI._0566_ vssd1 vssd1 vccd1 vccd1 AuI._0568_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4453_ MuI._0135_ MuI._0134_ vssd1 vssd1 vccd1 vccd1 MuI._0142_ sky130_fd_sc_hd__or2b_1
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05859_ _02907_ _04635_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__mux2_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4384_ MuI._3333_ MuI._3335_ vssd1 vssd1 vccd1 vccd1 MuI._0067_ sky130_fd_sc_hd__nor2_1
XFILLER_178_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0888__B1 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6123_ MuI._1963_ MuI._1964_ MuI._1976_ vssd1 vssd1 vccd1 vccd1 MuI._1979_ sky130_fd_sc_hd__and3_1
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6054_ MuI._3147_ MuI._1902_ vssd1 vssd1 vccd1 vccd1 MuI._1903_ sky130_fd_sc_hd__xor2_1
XANTENNA__12388__A2 _05233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _00772_ _00776_ _00777_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__and3_1
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5005_ MuI._0675_ MuI._0677_ vssd1 vssd1 vccd1 vccd1 MuI._0749_ sky130_fd_sc_hd__xor2_1
X_07111_ _06419_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[24\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_MuI._6176__A1 MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6176__B2 MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ _00707_ _00708_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13337__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4726__A2 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07042_ net28 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10634__B _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._792__A2 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5907_ MuI._1673_ MuI._1674_ vssd1 vssd1 vccd1 vccd1 MuI._1741_ sky130_fd_sc_hd__and2_1
XFILLER_88_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ _01605_ _01608_ _01609_ _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a211oi_2
XFILLER_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5838_ MuI._1651_ MuI._1664_ vssd1 vssd1 vccd1 vccd1 MuI._1665_ sky130_fd_sc_hd__xnor2_1
X_07944_ _00070_ _00071_ _00105_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__o21a_1
XFILLER_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._718_ AuI.pe._120_ AuI.pe._002_ AuI.pe._004_ AuI.pe._211_ AuI.pe._263_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._264_ sky130_fd_sc_hd__a221o_1
XFILLER_96_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5769_ MuI._1581_ MuI._1583_ MuI._1588_ vssd1 vssd1 vccd1 vccd1 MuI._1589_ sky130_fd_sc_hd__or3b_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07875_ _00485_ _00491_ _00492_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__nand3_1
XANTENNA__07662__C _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._649_ AuI.pe._125_ AuI.pe._078_ AuI.pe._119_ AuI.pe._071_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._199_ sky130_fd_sc_hd__a22o_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09614_ _02243_ _02244_ _02249_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__nand3_1
X_06826_ _03550_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__buf_4
XFILLER_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _02174_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__xor2_1
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06757_ _02808_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__and3_1
XANTENNA__08774__B _01387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ _02094_ _02095_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a21o_1
XFILLER_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11823__B2 _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ net2 _02064_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nor2_2
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08427_ _01038_ _01039_ _01042_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a21o_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10097__A _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._131_ FuI._015_ net137 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[2\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08358_ _00973_ _00974_ _00975_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__o21bai_1
XFILLER_196_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07309_ _06608_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__buf_6
XFILLER_192_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08289_ _00646_ _00647_ _00648_ _00649_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__and4_1
XFILLER_137_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ _03013_ _04983_ _03009_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__a22o_1
XANTENNA__13201__A _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _02559_ _02753_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or2_1
XFILLER_105_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__A2 _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _02970_ _04983_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__and2b_1
XFILLER_160_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1071__A3 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5142__A2 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09126__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1230_ AuI._0429_ AuI._0432_ vssd1 vssd1 vccd1 vccd1 AuI._0434_ sky130_fd_sc_hd__nor2_1
XANTENNA__07291__D _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ _05697_ _05701_ _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__or3_1
XAuI._1161_ AuI._0307_ AuI._0236_ AuI._0264_ vssd1 vssd1 vccd1 vccd1 AuI._0368_ sky130_fd_sc_hd__and3_1
XFILLER_90_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0814__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__A _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1092_ AuI._0254_ AuI._0300_ AuI._0301_ vssd1 vssd1 vccd1 vccd1 AuI._0303_ sky130_fd_sc_hd__and3_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _05626_ _05628_ _05540_ _05612_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a211oi_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _00878_ _05820_ _03444_ _00012_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a22o_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _05553_ _05554_ _05469_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__o21ai_2
XANTENNA_MuI._4414__A MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1348__C AuI._0542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4956__A2 MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ _04287_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__inv_2
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5229__B MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3675__D MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._501__A AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11567_ _03306_ _02790_ MuI.result\[9\] _02737_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4708__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13306_ _03134_ _06203_ _06204_ _06206_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__a311o_1
X_10518_ _06606_ _06601_ _05316_ _05380_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3972__B MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0945_ AuI._0150_ AuI._0156_ AuI._0096_ vssd1 vssd1 vccd1 vccd1 AuI._0157_ sky130_fd_sc_hd__a21o_1
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11498_ _04118_ _04120_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__nand2_1
XANTENNA__07747__C _00363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08205__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6810_ MuI._2731_ MuI._2733_ vssd1 vssd1 vccd1 vccd1 MuI._2734_ sky130_fd_sc_hd__or2b_1
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13237_ _03454_ _05595_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and2_1
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10449_ _03147_ _03148_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0876_ net112 net131 vssd1 vssd1 vccd1 vccd1 AuI._0096_ sky130_fd_sc_hd__xor2_1
XMuI._6741_ MuI._2474_ MuI._2467_ MuI._2471_ vssd1 vssd1 vccd1 vccd1 MuI._2658_ sky130_fd_sc_hd__and3_1
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3953_ MuI._3046_ MuI._3047_ MuI._3052_ vssd1 vssd1 vccd1 vccd1 MuI._3053_ sky130_fd_sc_hd__and3_1
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _03346_ _05467_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__nor2_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5133__A2 MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6672_ MuI._0282_ MuI._2581_ vssd1 vssd1 vccd1 vccd1 MuI._2582_ sky130_fd_sc_hd__nor2_1
X_12119_ _03658_ _04918_ _04818_ _04817_ _05047_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a32o_1
XMuI._3884_ MuI._2843_ MuI._2840_ MuI._2799_ MuI._2918_ vssd1 vssd1 vccd1 vccd1 MuI._2984_
+ sky130_fd_sc_hd__and4_1
X_13099_ _02632_ _05925_ _05998_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__a21o_1
XFILLER_111_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5623_ MuI._1400_ MuI._1410_ MuI._1427_ MuI._1376_ vssd1 vssd1 vccd1 vccd1 MuI._1429_
+ sky130_fd_sc_hd__or4b_1
XFILLER_78_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._503_ AuI.pe._059_ AuI.pe._049_ AuI.pe._063_ vssd1 vssd1 vccd1 vccd1 AuI.pe._064_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_38_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5554_ MuI._3403_ MuI._3245_ MuI._0020_ MuI._0304_ vssd1 vssd1 vccd1 vccd1 MuI._1353_
+ sky130_fd_sc_hd__and4_1
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1428_ AuI._0546_ AuI._0550_ vssd1 vssd1 vccd1 vccd1 AuI._0614_ sky130_fd_sc_hd__or2b_1
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07660_ net113 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._434_ AuI.pe._386_ AuI.pe._000_ AuI.pe._383_ AuI.pe._385_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._001_ sky130_fd_sc_hd__and4b_1
XFILLER_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4505_ MuI._0063_ MuI._0198_ vssd1 vssd1 vccd1 vccd1 MuI._0199_ sky130_fd_sc_hd__nand2_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5485_ MuI._2976_ MuI._0421_ MuI._1273_ MuI._1275_ vssd1 vssd1 vccd1 vccd1 MuI._1277_
+ sky130_fd_sc_hd__a211oi_1
XAuI._1359_ AuI._0552_ vssd1 vssd1 vccd1 vccd1 AuI._0553_ sky130_fd_sc_hd__inv_2
X_07591_ _00207_ _00208_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4519__A2_N MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4436_ MuI._0121_ MuI._0071_ MuI._3378_ MuI._0122_ vssd1 vssd1 vccd1 vccd1 MuI._0123_
+ sky130_fd_sc_hd__a211oi_1
X_09330_ _01912_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__nand2_1
XFILLER_179_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4367_ MuI._0035_ MuI._0036_ vssd1 vssd1 vccd1 vccd1 MuI._0048_ sky130_fd_sc_hd__nor2_1
X_09261_ _01876_ _01877_ _01669_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a21o_1
XFILLER_61_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6106_ MuI._1860_ MuI._1861_ vssd1 vssd1 vccd1 vccd1 MuI._1960_ sky130_fd_sc_hd__nor2_1
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6242__C MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ _00827_ _00828_ _00829_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__o21bai_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4298_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._3397_ vssd1 vssd1 vccd1
+ vccd1 MuI._3398_ sky130_fd_sc_hd__o31a_1
XFILLER_178_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09192_ _01798_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__or2_1
XMuI._6037_ MuI._3133_ MuI._3140_ vssd1 vssd1 vccd1 vccd1 MuI._1884_ sky130_fd_sc_hd__nand2_1
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10067__D _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ _00411_ _00413_ _00415_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07237__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B2 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout121_A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ _00460_ _00469_ _00468_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__a21o_1
XFILLER_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ net130 vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__buf_4
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B2 _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07954__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6857__C1 MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ _06488_ _04832_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__nand2_1
XFILLER_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07392__C _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _00536_ _00543_ _00544_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a21o_2
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12297__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1210__A0 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _00474_ _00475_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__nor2_1
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4218__B MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08000__D _00617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ net113 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__buf_4
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07789_ _00392_ _00393_ _00405_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__nand3_1
XFILLER_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09528_ _02153_ _02154_ _02156_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a21o_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _02066_ _02076_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__nor2_1
XFILLER_200_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08009__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10480__B1 _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ _05322_ _05323_ _05196_ _05199_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._5060__A1 MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5060__B2 MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._114_ FuI.a_operand\[26\] FuI._037_ FuI._054_ vssd1 vssd1 vccd1 vccd1 FuI._026_
+ sky130_fd_sc_hd__or3_1
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04193_ _04194_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI._1277__A0 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__A2 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ _04119_ _04120_ _04116_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a21o_1
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _02991_ _02989_ _02990_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._5065__A MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ _04028_ _04045_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__nand3_2
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07286__D _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ _05915_ _05916_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__nand2_1
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10234_ _03626_ _05788_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__and2b_1
XANTENNA_input51_A b_operand[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12797__A1_N _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07400__A1 _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10165_ _00566_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor2_2
XFILLER_94_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13485__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _02715_ _02714_ _02753_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__and3_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1213_ AuI._0416_ AuI._0417_ vssd1 vssd1 vccd1 vccd1 AuI._0418_ sky130_fd_sc_hd__or2_2
XFILLER_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5270_ MuI.a_operand\[14\] MuI._3402_ MuI._3396_ MuI.a_operand\[15\] vssd1 vssd1
+ vccd1 vccd1 MuI._1040_ sky130_fd_sc_hd__a22oi_2
X_12806_ _05685_ _02904_ _02926_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__mux2_1
XAuI._1144_ AuI._0274_ AuI._0312_ vssd1 vssd1 vccd1 vccd1 AuI._0352_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3967__B MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10998_ _03738_ _03739_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or2_1
XMuI._4221_ MuI._3315_ MuI._3320_ vssd1 vssd1 vccd1 vccd1 MuI._3321_ sky130_fd_sc_hd__and2_1
XANTENNA__11819__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _05451_ _05453_ _05540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08664__B1 _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1075_ AuI._0283_ AuI._0285_ AuI._0208_ vssd1 vssd1 vccd1 vccd1 AuI._0286_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4152_ MuI._3250_ MuI._3251_ vssd1 vssd1 vccd1 vccd1 MuI._3252_ sky130_fd_sc_hd__nand2_1
XFILLER_148_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ _05535_ _05536_ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__a21o_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4083_ MuI._2870_ MuI._2877_ MuI._2872_ vssd1 vssd1 vccd1 vccd1 MuI._3183_ sky130_fd_sc_hd__o21ai_1
XFILLER_191_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _04406_ _04407_ _04408_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o21ai_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ _05289_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__or3_1
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5354__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__B _02637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0928_ net5 net37 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0140_ sky130_fd_sc_hd__mux2_1
XFILLER_125_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4985_ MuI._0746_ MuI._1164_ MuI._0245_ MuI._0321_ vssd1 vssd1 vccd1 vccd1 MuI._0727_
+ sky130_fd_sc_hd__and4_1
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._0859_ net122 AuI._0074_ AuI._0078_ net6 vssd1 vssd1 vccd1 vccd1 AuI._0079_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_98_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6724_ MuI._2637_ MuI._2639_ vssd1 vssd1 vccd1 vccd1 MuI._2640_ sky130_fd_sc_hd__nor2_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5106__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3936_ MuI._2787_ MuI._2407_ MuI._3022_ MuI._3023_ vssd1 vssd1 vccd1 vccd1 MuI._3036_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08830_ _01441_ _01446_ _01445_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a21o_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6655_ MuI._2553_ MuI._2555_ MuI._1442_ vssd1 vssd1 vccd1 vccd1 MuI._2564_ sky130_fd_sc_hd__or3b_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3867_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._2967_ sky130_fd_sc_hd__clkbuf_4
X_08761_ _01373_ _01378_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__and2_1
XFILLER_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5606_ MuI._1398_ MuI._1399_ MuI._1393_ MuI._1397_ vssd1 vssd1 vccd1 vccd1 MuI._1410_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07712_ _00285_ _00296_ vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__and2b_1
XMuI._6586_ MuI._0295_ MuI._0317_ MuI._2487_ MuI.a_operand\[23\] vssd1 vssd1 vccd1
+ vccd1 MuI._2488_ sky130_fd_sc_hd__a211o_1
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3798_ MuI._2871_ vssd1 vssd1 vccd1 vccd1 MuI._2898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08692_ _01066_ _01067_ _01117_ _01118_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__and4_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5537_ MuI._1330_ MuI._1333_ vssd1 vssd1 vccd1 vccd1 MuI._1334_ sky130_fd_sc_hd__or2b_1
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07643_ _00257_ _00260_ vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__nor2_1
XFILLER_199_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._417_ AuI.pe._383_ vssd1 vssd1 vccd1 vccd1 AuI.pe._384_ sky130_fd_sc_hd__clkbuf_2
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5468_ MuI._1250_ MuI._1251_ MuI._1256_ vssd1 vssd1 vccd1 vccd1 MuI._1258_ sky130_fd_sc_hd__nand3_1
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07574_ _00189_ _00190_ _00191_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__or3_1
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09447__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__B _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4419_ MuI._0099_ MuI._0102_ MuI._0103_ vssd1 vssd1 vccd1 vccd1 MuI._0104_ sky130_fd_sc_hd__o21ba_1
X_09313_ net111 _00030_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__nand2_1
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07014__A _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5399_ MuI._1181_ vssd1 vssd1 vccd1 vccd1 MuI._1182_ sky130_fd_sc_hd__inv_2
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3840__A2 MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09244_ _01650_ _01857_ _01860_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a211oi_2
XFILLER_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06853__A _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ _01791_ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10375__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09586__D _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08126_ _00725_ _00726_ _00743_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__o21ba_1
XFILLER_181_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__B _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08057_ _00505_ _00513_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__or2b_1
XFILLER_162_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12506__A2 _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ _05509_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_162_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08959_ _01575_ _01568_ _01569_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nand3_1
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _00299_ _00231_ _00530_ _06666_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and4_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10921_ _03509_ _03510_ _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__a21o_1
XFILLER_17_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _03579_ _03580_ _03581_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a21o_1
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08665__D net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10269__B _00708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10783_ _03482_ _03479_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or2b_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3831__A2 MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12522_ _05379_ _02850_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__nor2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nand2_1
XFILLER_173_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11404_ _02773_ _04178_ _02750_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__o21ai_1
XANTENNA_MuI._5507__B MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09071__B1 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12384_ _05230_ _05231_ _05120_ _05122_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__a211o_1
XFILLER_181_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09610__A2 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _03525_ _04531_ _03866_ _03865_ _04660_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a32o_2
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11266_ _00878_ _05649_ _03449_ _00877_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a22oi_1
XFILLER_180_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11705__B1 _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4770_ MuI._0465_ MuI._0473_ MuI._0475_ vssd1 vssd1 vccd1 vccd1 MuI._0490_ sky130_fd_sc_hd__nand3_1
X_10217_ _02899_ _02865_ _02863_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
X_13005_ _05897_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__xor2_2
XFILLER_140_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11197_ _03745_ _03747_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__nand2_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3721_ MuI._2813_ MuI._2786_ MuI._2363_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._2821_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4784__D MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _02814_ _02817_ _02822_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or4_2
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6440_ MuI._2282_ MuI._2310_ MuI._2318_ vssd1 vssd1 vccd1 vccd1 MuI._2327_ sky130_fd_sc_hd__o21ai_1
XFILLER_208_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3652_ MuI._2429_ vssd1 vssd1 vccd1 vccd1 MuI._2528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_208_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ _02750_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__buf_6
XANTENNA__06938__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6371_ MuI._2250_ vssd1 vssd1 vccd1 vccd1 MuI._2251_ sky130_fd_sc_hd__inv_2
XMuI._3583_ MuI._1340_ MuI._1527_ vssd1 vssd1 vccd1 vccd1 MuI._1769_ sky130_fd_sc_hd__or2_1
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5322_ MuI._1091_ MuI._1092_ MuI._1096_ vssd1 vssd1 vccd1 vccd1 MuI._1097_ sky130_fd_sc_hd__a21o_1
XFuI._134__140 vssd1 vssd1 vccd1 vccd1 FuI._134__140/HI net140 sky130_fd_sc_hd__conb_1
XFILLER_63_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12992__B1_N _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5253_ MuI._1018_ MuI._1019_ MuI._1020_ vssd1 vssd1 vccd1 vccd1 MuI._1022_ sky130_fd_sc_hd__nand3b_1
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1127_ AuI._0206_ AuI._0192_ AuI._0264_ vssd1 vssd1 vccd1 vccd1 AuI._0336_ sky130_fd_sc_hd__and3_1
XMuI._4204_ MuI._3302_ MuI._3303_ vssd1 vssd1 vccd1 vccd1 MuI._3304_ sky130_fd_sc_hd__nor2b_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5184_ MuI._0939_ MuI._0945_ vssd1 vssd1 vccd1 vccd1 MuI._0946_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12984__A2 _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ _06580_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__buf_4
XAuI._1058_ AuI._0164_ AuI._0169_ AuI._0214_ vssd1 vssd1 vccd1 vccd1 AuI._0269_ sky130_fd_sc_hd__and3_1
XFILLER_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4135_ MuI._0878_ MuI._2385_ MuI._2820_ MuI._2821_ vssd1 vssd1 vccd1 vccd1 MuI._3235_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10195__A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12197__B1 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07919__D _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4066_ MuI._3073_ MuI._3074_ MuI._3072_ vssd1 vssd1 vccd1 vccd1 MuI._3166_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4783__B1 MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4321__B MuI._3420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _02588_ _02590_ _02591_ _02034_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a211oi_2
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4968_ MuI._0632_ MuI._0634_ MuI._0645_ vssd1 vssd1 vccd1 vccd1 MuI._0708_ sky130_fd_sc_hd__a21oi_1
X_09862_ _02490_ _02491_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__and3_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08112__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3919_ MuI._2938_ MuI._3012_ MuI._3017_ vssd1 vssd1 vccd1 vccd1 MuI._3019_ sky130_fd_sc_hd__or3_1
XMuI._6707_ MuI._2608_ MuI._2612_ MuI._2617_ MuI._2620_ vssd1 vssd1 vccd1 vccd1 MuI._2621_
+ sky130_fd_sc_hd__nor4_1
XFILLER_140_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5152__B MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ _01423_ _01429_ _01430_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a21o_1
XANTENNA__07009__A _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4899_ MuI._0621_ MuI._0629_ MuI._0631_ vssd1 vssd1 vccd1 vccd1 MuI._0632_ sky130_fd_sc_hd__a21o_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _02347_ _02443_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__nor2_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6638_ MuI._1438_ MuI._1442_ vssd1 vssd1 vccd1 vccd1 MuI._2545_ sky130_fd_sc_hd__nor2_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _02840_ _04251_ _01359_ _01360_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4991__B MuI._0726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06848__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6569_ MuI._2464_ MuI._2458_ MuI._2456_ vssd1 vssd1 vccd1 vccd1 MuI._2469_ sky130_fd_sc_hd__o21a_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07670__C _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _01225_ _01224_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__and2b_1
XFILLER_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11192__C _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07626_ _00240_ _00241_ _00242_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__a21o_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5263__A1 MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__B _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07557_ net106 _06476_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__nand2_1
XANTENNA__12424__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__B _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12424__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07488_ _00070_ _00071_ _00105_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__or3_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09840__A2 _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _01677_ _01678_ _01766_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__or3_1
XFILLER_195_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07829__D _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ net107 net66 _00082_ net36 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__and4_1
XFILLER_107_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _00231_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__buf_4
X_09089_ _01680_ _01695_ _01694_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a21o_1
XANTENNA__12524__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__xor2_4
XFILLER_190_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08303__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09356__A1 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09356__B2 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _03794_ _03795_ _03780_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a21o_1
XFILLER_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _02650_ _02653_ _02654_ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__or3_1
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3798__A MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input14_A a_operand[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _02808_ _02851_ _05895_ _05970_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__nand4_2
XANTENNA_MuI._6174__A MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ _03636_ _03638_ _03596_ _03597_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a211oi_1
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ _04693_ _04675_ _04676_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nand3_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10835_ _03559_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nand3_1
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6203__B1 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ _02768_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A1 _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10977__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _02865_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__inv_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13485_ MuI.result\[31\] _02739_ _02938_ AuI.result\[31\] _06400_ vssd1 vssd1 vccd1
+ vccd1 _06401_ sky130_fd_sc_hd__a221o_1
X_10697_ _03234_ _03236_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__nand2_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12179__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5237__B MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ _05267_ _05174_ _05287_ _05288_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__o211ai_4
XFILLER_173_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5940_ MuI._1775_ MuI._1749_ MuI._1776_ MuI._0733_ vssd1 vssd1 vccd1 vccd1 MuI._1777_
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12367_ _03744_ _04983_ _05085_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__a31o_1
XAuI.pe._820_ AuI.pe._330_ AuI.pe._341_ AuI.pe._339_ vssd1 vssd1 vccd1 vccd1 AuI.pe._359_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_114_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5871_ MuI._1682_ MuI._1683_ MuI._1698_ MuI._1699_ vssd1 vssd1 vccd1 vccd1 MuI._1701_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_154_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output82_A net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11318_ _04067_ _04069_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a21oi_2
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12298_ _02795_ _05017_ _02792_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o21bai_1
XAuI.pe._751_ AuI.pe.significand\[22\] AuI.pe._291_ AuI.pe._294_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._295_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10462__B _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4822_ MuI._0419_ MuI._0546_ vssd1 vssd1 vccd1 vccd1 MuI._0547_ sky130_fd_sc_hd__nor2_1
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11249_ _02129_ _01988_ _04011_ _02756_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o211a_1
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._682_ AuI.pe._084_ AuI.pe._133_ AuI.pe._228_ AuI.pe._229_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._230_ sky130_fd_sc_hd__a211o_1
XANTENNA__09898__A2 _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4753_ MuI._0465_ MuI._0470_ vssd1 vssd1 vccd1 vccd1 MuI._0472_ sky130_fd_sc_hd__and2_1
XFILLER_121_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3704_ MuI._2802_ MuI._2803_ MuI._2671_ MuI._2528_ vssd1 vssd1 vccd1 vccd1 MuI._2804_
+ sky130_fd_sc_hd__and4_1
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4684_ MuI._0392_ MuI._0393_ MuI._0395_ vssd1 vssd1 vccd1 vccd1 MuI._0396_ sky130_fd_sc_hd__a21bo_1
X_06790_ _03163_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__clkbuf_8
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6423_ MuI._2303_ MuI._2301_ vssd1 vssd1 vccd1 vccd1 MuI._2309_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3635_ MuI.a_operand\[8\] vssd1 vssd1 vccd1 vccd1 MuI._2341_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08586__C _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6354_ MuI._2207_ MuI._2230_ vssd1 vssd1 vccd1 vccd1 MuI._2233_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._3501__A MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3566_ MuI._1109_ MuI._1252_ MuI._1571_ vssd1 vssd1 vccd1 vccd1 MuI._1582_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10665__B1 _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _01070_ _01076_ _01075_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__a21o_1
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5305_ MuI._1074_ MuI._1078_ vssd1 vssd1 vccd1 vccd1 MuI._1079_ sky130_fd_sc_hd__nor2_1
XANTENNA_AuI.pe._638__A1 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07411_ net44 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__buf_4
XFILLER_196_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6285_ MuI._2119_ MuI._2125_ MuI._2117_ vssd1 vssd1 vccd1 vccd1 MuI._2157_ sky130_fd_sc_hd__a21oi_1
XMuI._3497_ MuI._0350_ MuI._0636_ MuI._0592_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._0823_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12406__A1 AuI.result\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ _00993_ _00996_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__and2b_1
XANTENNA__12406__B2 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5236_ MuI._2583_ MuI._0315_ vssd1 vssd1 vccd1 vccd1 MuI._1003_ sky130_fd_sc_hd__nand2_1
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07342_ _02107_ _06495_ net129 net128 vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__and4_1
XFILLER_176_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10130__A_N _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5167_ MuI._0924_ MuI._0925_ MuI._0905_ vssd1 vssd1 vccd1 vccd1 MuI._0927_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _06556_ _06557_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._3874__C MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4118_ MuI._2704_ MuI._2803_ MuI._2528_ MuI._2539_ vssd1 vssd1 vccd1 vccd1 MuI._3218_
+ sky130_fd_sc_hd__and4_1
X_09012_ _01291_ _01292_ _01294_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and3_1
XFILLER_192_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5098_ MuI._0848_ MuI._0849_ MuI._0850_ vssd1 vssd1 vccd1 vccd1 MuI._0851_ sky130_fd_sc_hd__or3_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4049_ MuI._3147_ MuI._3148_ vssd1 vssd1 vccd1 vccd1 MuI._3149_ sky130_fd_sc_hd__nand2_1
XFILLER_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11393__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6259__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5181__B1 MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _02484_ _02486_ _02520_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__and3_1
XANTENNA__13134__A2 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _02498_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__xnor2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A a_operand[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5633__A2_N MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _02229_ net115 _06437_ _02442_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22oi_1
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ net18 vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__clkbuf_4
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5610__B MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ _02550_ _04531_ _01343_ _01344_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__a31o_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12645__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12645__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _01135_ _01136_ _01173_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__or3_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4226__B MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._629__B2 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12504__A1_N _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07609_ _00116_ _00117_ _00115_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__a21bo_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08520__A_N _01102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ _01206_ _06446_ _00303_ _00921_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a22o_1
XFILLER_168_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13204__A _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _03178_ _03140_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or2b_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07202__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ _00162_ _03082_ _00789_ _00164_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a22o_1
XANTENNA__11620__A2 _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4242__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__D _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _00058_ _00421_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__nand2_4
X_13270_ _06167_ _06116_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12762__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11659__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ _03163_ _03425_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__nand2_1
XFILLER_170_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _04939_ _04981_ _04982_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3_1
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10282__B _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _03851_ _03853_ _02925_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__mux2_1
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1530_ AuI._0710_ AuI._0713_ vssd1 vssd1 vccd1 vccd1 AuI._0714_ sky130_fd_sc_hd__nand2_1
XFILLER_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12083_ _02894_ _00046_ _00783_ _05884_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and4_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11034_ _03621_ _03629_ _03628_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07872__A _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1461_ AuI._0358_ AuI._0361_ vssd1 vssd1 vccd1 vccd1 AuI._0647_ sky130_fd_sc_hd__and2b_1
XFILLER_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12884__B2 _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11394__A _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1392_ AuI._0580_ AuI._0582_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[21\]
+ sky130_fd_sc_hd__xnor2_4
XFILLER_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3486__B1 MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12985_ _05875_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__xor2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__A2 _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _04749_ _04750_ _04554_ _04598_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211oi_2
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._504__A AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _00124_ _05316_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__nand2_2
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6070_ MuI._1872_ MuI._1877_ MuI._1870_ vssd1 vssd1 vccd1 vccd1 MuI._1920_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10818_ _03543_ _03544_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
XFILLER_159_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5021_ MuI._0611_ MuI._0764_ MuI._0763_ MuI._0760_ vssd1 vssd1 vccd1 vccd1 MuI._0766_
+ sky130_fd_sc_hd__a211o_1
X_11798_ _04600_ _04601_ _04469_ _04471_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07112__A _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10749_ _03219_ _03275_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13468_ _06370_ _06371_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06951__A _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09477__A2_N _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__B _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _01146_ _03425_ _03449_ _01147_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a22oi_1
XFILLER_173_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _03314_ _06305_ _06306_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__a31o_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5923_ MuI._1756_ MuI._1757_ vssd1 vssd1 vccd1 vccd1 MuI._1759_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._803_ AuI.pe._273_ AuI.pe._375_ AuI.pe._049_ vssd1 vssd1 vccd1 vccd1 AuI.pe._342_
+ sky130_fd_sc_hd__nor3_1
XMuI._5854_ MuI._1679_ MuI._1680_ MuI._1581_ MuI._1668_ vssd1 vssd1 vccd1 vccd1 MuI._1683_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _00052_ _00054_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__xnor2_1
XMuI._4805_ MuI._0523_ MuI._0528_ vssd1 vssd1 vccd1 vccd1 MuI._0529_ sky130_fd_sc_hd__nor2_1
XAuI.pe._734_ AuI.pe._046_ AuI.pe._225_ AuI.pe._277_ AuI.pe._084_ AuI.pe._278_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._279_ sky130_fd_sc_hd__a221o_1
XMuI._5785_ MuI._1605_ MuI._1606_ vssd1 vssd1 vccd1 vccd1 MuI._1607_ sky130_fd_sc_hd__xnor2_1
X_06911_ _02151_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__clkbuf_2
XAuI._1659_ AuI.exponent_sub\[4\] AuI._0599_ AuI._0698_ vssd1 vssd1 vccd1 vccd1 AuI._0013_
+ sky130_fd_sc_hd__o21a_1
XFILLER_68_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07891_ _00507_ _00508_ _06439_ _06443_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__and4bb_1
XAuI.pe._665_ AuI.pe._033_ AuI.pe._397_ AuI.pe._213_ AuI.pe._014_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._214_ sky130_fd_sc_hd__a22o_1
XANTENNA__08597__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__B _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4736_ MuI._0451_ MuI._0452_ vssd1 vssd1 vccd1 vccd1 MuI._0453_ sky130_fd_sc_hd__or2_1
X_09630_ _02265_ _02266_ _02237_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06842_ _03722_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__C _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._596_ AuI.pe._149_ AuI.pe._379_ vssd1 vssd1 vccd1 vccd1 AuI.pe._150_ sky130_fd_sc_hd__nor2_4
XMuI._4667_ MuI.a_operand\[19\] MuI._0017_ MuI._0018_ MuI.a_operand\[20\] vssd1 vssd1
+ vccd1 vccd1 MuI._0377_ sky130_fd_sc_hd__a22oi_1
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4972__D MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ _02981_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[16\] sky130_fd_sc_hd__clkbuf_1
X_09561_ _02191_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__xnor2_1
XMuI._6406_ MuI._2285_ MuI._2278_ MuI._2288_ vssd1 vssd1 vccd1 vccd1 MuI._2290_ sky130_fd_sc_hd__nand3_1
XMuI._3618_ MuI._1417_ MuI._1516_ vssd1 vssd1 vccd1 vccd1 MuI._2154_ sky130_fd_sc_hd__or2b_1
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08512_ _01128_ _01127_ _01062_ _01060_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__o211a_1
XMuI._4598_ MuI._0291_ MuI._0299_ MuI._0300_ vssd1 vssd1 vccd1 vccd1 MuI._0301_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09492_ _02110_ _02111_ _02116_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a21o_1
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6337_ MuI._0889_ MuI._1043_ MuI._1945_ vssd1 vssd1 vccd1 vccd1 MuI._2214_ sky130_fd_sc_hd__a21oi_1
XANTENNA_AuI.pe._414__A AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3549_ MuI._0581_ MuI._1164_ MuI._0757_ vssd1 vssd1 vccd1 vccd1 MuI._1395_ sky130_fd_sc_hd__and3_1
XFILLER_51_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ _01057_ _01058_ _01059_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__nand3_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6268_ MuI._2018_ MuI._2026_ vssd1 vssd1 vccd1 vccd1 MuI._2138_ sky130_fd_sc_hd__and2_1
XANTENNA__08059__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _00988_ _00991_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__or2b_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08118__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5219_ MuI._0847_ MuI._0982_ MuI._0983_ vssd1 vssd1 vccd1 vccd1 MuI._0984_ sky130_fd_sc_hd__a21bo_1
XFILLER_177_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ _06624_ _06625_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__and2b_1
XANTENNA__07022__A _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6199_ MuI._2056_ MuI._2061_ vssd1 vssd1 vccd1 vccd1 MuI._2062_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07806__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4062__A MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07806__B2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07256_ _06553_ _06555_ _06554_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._6194__A2 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6688__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06861__A _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13355__A2 _06261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07187_ net111 vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__buf_4
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12563__B1 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12315__B1 _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07692__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12072__B_N _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09828_ _02477_ _02479_ _02438_ _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a211oi_2
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07742__B1 _00359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09759_ _02364_ _02355_ _02363_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nand3_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05629_ _05630_ _05645_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__o21ba_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _04516_ _04517_ _04513_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__a21o_1
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__xnor2_4
XFILLER_168_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _03314_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__buf_4
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _04225_ _04226_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__a21o_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4403__C MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ _06231_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__nor2_1
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ _03238_ _03240_ _03220_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0961_ AuI._0164_ AuI._0169_ AuI._0172_ vssd1 vssd1 vccd1 vccd1 AuI._0173_ sky130_fd_sc_hd__and3_1
XFILLER_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06771__A _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ _02833_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or2_1
X_10465_ _02985_ _02988_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nand2_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10293__A _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0892_ net129 vssd1 vssd1 vccd1 vccd1 AuI._0112_ sky130_fd_sc_hd__inv_2
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12204_ _02959_ _03444_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__nand2_1
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13184_ _02645_ _06089_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__o21a_1
XFILLER_108_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10396_ _00788_ _00794_ _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a21oi_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _04959_ _04963_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__nand3_1
XANTENNA__08773__A2 _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5696__A1 MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1513_ AuI._0698_ vssd1 vssd1 vccd1 vccd1 AuI._0699_ sky130_fd_sc_hd__buf_2
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _04881_ _04882_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__o21ai_2
XMuI._5570_ MuI._1365_ MuI._1367_ MuI._1368_ MuI._1369_ vssd1 vssd1 vccd1 vccd1 MuI._1370_
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__09722__A1 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__B2 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1444_ AuI._0503_ AuI._0493_ vssd1 vssd1 vccd1 vccd1 AuI._0630_ sky130_fd_sc_hd__nor2_1
X_11017_ _03759_ _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10868__B1 _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._450_ AuI.pe.significand\[7\] AuI.pe._370_ AuI.pe._374_ AuI.pe.significand\[6\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._017_ sky130_fd_sc_hd__or4b_1
XMuI._4521_ MuI._3000_ MuI._1791_ MuI._0088_ MuI._3362_ vssd1 vssd1 vccd1 vccd1 MuI._0216_
+ sky130_fd_sc_hd__and4_1
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5250__B MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1375_ AuI._0257_ AuI._0565_ AuI._0566_ vssd1 vssd1 vccd1 vccd1 AuI._0567_ sky130_fd_sc_hd__and3_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4147__A MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4452_ MuI._0138_ MuI._0016_ vssd1 vssd1 vccd1 vccd1 MuI._0140_ sky130_fd_sc_hd__xor2_1
XFILLER_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _02805_ _02809_ _05685_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a31oi_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06946__A _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4383_ MuI._0041_ MuI._0046_ vssd1 vssd1 vccd1 vccd1 MuI._0066_ sky130_fd_sc_hd__or2b_1
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11919_ _04730_ _04731_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a21o_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6122_ MuI._1963_ MuI._1964_ MuI._1976_ vssd1 vssd1 vccd1 vccd1 MuI._1977_ sky130_fd_sc_hd__a21oi_1
X_12899_ _05710_ _05711_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__and2b_1
XFILLER_60_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6053_ MuI._1885_ MuI._1900_ vssd1 vssd1 vccd1 vccd1 MuI._1902_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5004_ MuI._0555_ MuI._0745_ MuI._0744_ vssd1 vssd1 vccd1 vccd1 MuI._0748_ sky130_fd_sc_hd__a21o_1
XFILLER_186_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07110_ _05531_ _06414_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and2_1
XFILLER_186_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _00495_ _00497_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__nor2_2
XFILLER_174_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07041_ _05863_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[29\] sky130_fd_sc_hd__clkbuf_2
XANTENNA__13337__A2 _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5906_ MuI._1738_ MuI._1739_ vssd1 vssd1 vccd1 vccd1 MuI._1740_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12622__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _01470_ _01471_ _01480_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5837_ MuI._1652_ MuI._1663_ vssd1 vssd1 vccd1 vccd1 MuI._1664_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._409__A AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__A1_N _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07943_ _00553_ _00559_ _00545_ _00560_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__o211ai_4
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08401__A _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._717_ AuI.pe._386_ AuI.pe._006_ AuI.pe._040_ AuI.pe._385_ AuI.pe._262_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._263_ sky130_fd_sc_hd__a221o_1
XMuI._5768_ MuI._1584_ MuI._1587_ vssd1 vssd1 vccd1 vccd1 MuI._1588_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07874_ _00489_ _00490_ _00486_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a21o_1
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__D _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._648_ AuI.pe._030_ AuI.pe._084_ AuI.pe._197_ AuI.pe._150_ AuI.pe._059_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._198_ sky130_fd_sc_hd__a32o_1
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4719_ MuI._0294_ MuI._0428_ vssd1 vssd1 vccd1 vccd1 MuI._0434_ sky130_fd_sc_hd__nor2_1
X_09613_ _02243_ _02244_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a21o_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5699_ MuI._1506_ MuI._1510_ MuI._1511_ vssd1 vssd1 vccd1 vccd1 MuI._1512_ sky130_fd_sc_hd__and3_1
X_06825_ _03539_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._579_ AuI.pe._378_ AuI.pe._026_ AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 AuI.pe._134_
+ sky130_fd_sc_hd__a21o_1
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11762__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _02057_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__and2b_1
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06756_ _02797_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__buf_8
XANTENNA__06856__A _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ net1 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__buf_2
X_09475_ _02097_ _02098_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o21bai_1
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _00992_ _01000_ _00999_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a21o_1
XFuI._130_ FuI._014_ net136 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[1\] sky130_fd_sc_hd__dlxtn_1
XFILLER_200_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _06494_ _06495_ _05241_ _05305_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__and4_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__B _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07308_ _06600_ _06607_ _06608_ _04789_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and4bb_1
XFILLER_165_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ _00646_ _00647_ _00648_ _00649_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__a22oi_2
XFILLER_109_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07239_ _06462_ _06464_ _06459_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13201__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10250_ _02559_ _02753_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nand2_1
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__inv_2
XANTENNA_MuI._4259__A1_N MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5678__A1 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4350__A1 MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4350__B2 MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09126__B _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ _05700_ _05698_ _05699_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor3_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1160_ AuI._0304_ AuI._0320_ AuI._0342_ AuI._0358_ vssd1 vssd1 vccd1 vccd1 AuI._0367_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__06766__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12487__B _05341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1091_ AuI._0300_ AuI._0301_ AuI._0254_ vssd1 vssd1 vccd1 vccd1 AuI._0302_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ _05540_ _05612_ _05626_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__o211a_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11704_ _00877_ _00878_ _05820_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__and3_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4405__A2 MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ _05469_ _05553_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__or3_4
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4414__B MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11635_ _04424_ _04425_ _04365_ _04249_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__a211o_1
XFILLER_168_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0830__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11566_ _02604_ _04542_ _02744_ _02945_ _04467_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__a32o_1
XANTENNA__09640__B1 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _03314_ _06208_ _06209_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a31o_1
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ _02808_ _03047_ _06477_ _02765_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a22oi_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0944_ AuI._0155_ AuI._0097_ vssd1 vssd1 vccd1 vccd1 AuI._0156_ sky130_fd_sc_hd__or2b_1
XANTENNA_AuI._1364__C AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _04276_ _04277_ _04272_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21o_1
XANTENNA__08205__B _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ MuI.result\[25\] _02738_ _04642_ _05531_ _06144_ vssd1 vssd1 vccd1 vccd1
+ _06145_ sky130_fd_sc_hd__a221o_1
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0875_ AuI._0046_ AuI._0093_ AuI._0028_ AuI._0094_ vssd1 vssd1 vccd1 vccd1 AuI._0095_
+ sky130_fd_sc_hd__o211ai_1
X_10448_ _02962_ _02966_ _02963_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o21ba_1
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3952_ MuI._3048_ MuI._3051_ vssd1 vssd1 vccd1 vccd1 MuI._3052_ sky130_fd_sc_hd__xnor2_1
XMuI._6740_ MuI._2652_ vssd1 vssd1 vccd1 vccd1 MuI._2657_ sky130_fd_sc_hd__clkinv_2
XANTENNA__11847__A _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13167_ _06063_ _06071_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__or2_1
X_10379_ _02539_ _03071_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__nand4_1
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6671_ MuI._1836_ MuI._1840_ MuI._0786_ vssd1 vssd1 vccd1 vccd1 MuI._2581_ sky130_fd_sc_hd__o21ba_1
XMuI._3883_ MuI.b_operand\[14\] MuI._2616_ vssd1 vssd1 vccd1 vccd1 MuI._2983_ sky130_fd_sc_hd__nand2_1
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12118_ _04945_ _04946_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__xor2_1
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _02632_ _05998_ _05925_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nand3_2
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5622_ MuI._1413_ MuI._1426_ vssd1 vssd1 vccd1 vccd1 MuI._1427_ sky130_fd_sc_hd__nand2_1
XFILLER_78_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12049_ _04614_ _04615_ _04761_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__nor3_1
XAuI.pe._502_ AuI.pe._062_ vssd1 vssd1 vccd1 vccd1 AuI.pe._063_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5553_ MuI._0228_ MuI._3397_ MuI._0305_ MuI._3403_ vssd1 vssd1 vccd1 vccd1 MuI._1352_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1427_ AuI._0560_ AuI._0557_ vssd1 vssd1 vccd1 vccd1 AuI._0613_ sky130_fd_sc_hd__and2b_1
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4504_ MuI._0060_ MuI._0062_ vssd1 vssd1 vccd1 vccd1 MuI._0198_ sky130_fd_sc_hd__or2_1
XAuI.pe._433_ AuI.pe.significand\[20\] vssd1 vssd1 vccd1 vccd1 AuI.pe._000_ sky130_fd_sc_hd__inv_2
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5484_ MuI._1273_ MuI._1275_ MuI._2976_ MuI._0420_ vssd1 vssd1 vccd1 vccd1 MuI._1276_
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1358_ AuI._0526_ AuI._0527_ AuI._0544_ AuI._0543_ vssd1 vssd1 vccd1 vccd1 AuI._0552_
+ sky130_fd_sc_hd__a31oi_1
X_07590_ _00204_ _00206_ _00205_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a21o_1
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4644__A2 MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4435_ MuI._3357_ MuI._3358_ MuI._3377_ vssd1 vssd1 vccd1 vccd1 MuI._0122_ sky130_fd_sc_hd__o21a_1
XANTENNA__12397__B _02584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11266__B1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__A _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1289_ AuI._0263_ AuI._0371_ vssd1 vssd1 vccd1 vccd1 AuI._0488_ sky130_fd_sc_hd__nor2_1
XFILLER_206_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4605__A MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4366_ MuI._0041_ MuI._0046_ vssd1 vssd1 vccd1 vccd1 MuI._0047_ sky130_fd_sc_hd__xnor2_2
X_09260_ _01669_ _01876_ _01877_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nand3_2
XMuI._6105_ MuI._1860_ MuI._1861_ vssd1 vssd1 vccd1 vccd1 MuI._1959_ sky130_fd_sc_hd__and2_1
XFILLER_178_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11018__B1 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _06469_ _02194_ net19 net20 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__and4_1
XMuI._4297_ MuI._3396_ vssd1 vssd1 vccd1 vccd1 MuI._3397_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._6242__D MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _01798_ _01799_ _01807_ _01808_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__nor4_1
XFILLER_193_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10926__A _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6036_ MuI._1881_ MuI._1882_ vssd1 vssd1 vccd1 vccd1 MuI._1883_ sky130_fd_sc_hd__xnor2_1
X_08142_ _00756_ _00757_ _00758_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__o21ai_1
XFILLER_193_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07237__A2 _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _00689_ _00690_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__xnor2_4
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4340__A MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__B1 _05376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07024_ _05682_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[26\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_MuI._5155__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__A2 _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__B _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6857__B1 MuI._2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6869_ MuI._2497_ MuI._0240_ vssd1 vssd1 vccd1 vccd1 MuI._2770_ sky130_fd_sc_hd__and2b_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08975_ _01459_ _01458_ _01457_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21o_1
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07926_ _06597_ _06615_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ _00472_ _00473_ _00204_ _00207_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__o211a_1
XFILLER_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1210__A1 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4218__C MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _03357_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[23\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07788_ _00392_ _00393_ _00405_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a21o_1
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09527_ _02153_ _02154_ _02156_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nand3_1
X_06739_ _02604_ _02615_ _02162_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__and3_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4515__A MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _02765_ _03895_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10480__A1 _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08009__C _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08409_ _01022_ _01023_ _01026_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__nand3_1
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10480__B2 _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._113_ FuI._023_ FuI._061_ FuI._054_ vssd1 vssd1 vccd1 vccd1 FuI._025_ sky130_fd_sc_hd__or3_1
X_09389_ _02005_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _04058_ _04060_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__nand2_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1277__A1 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5346__A MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _04116_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nand3_2
XFILLER_153_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ _02989_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5065__B MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11282_ _04043_ _04044_ _03916_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a21o_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4571__A1 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _05864_ _05832_ _05914_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nand3_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10233_ _02917_ _05917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__and2_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0809__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input44_A b_operand[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _02765_ _04736_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__nor2_1
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5520__B1 MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10095_ _02767_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__and2_1
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08976__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08361__B1 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1212_ AuI._0412_ AuI._0414_ AuI._0415_ vssd1 vssd1 vccd1 vccd1 AuI._0417_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0960__A0 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _02866_ _05594_ _02867_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__o21ba_1
XAuI._1143_ AuI._0263_ AuI._0350_ vssd1 vssd1 vccd1 vccd1 AuI._0351_ sky130_fd_sc_hd__nand2_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4220_ MuI._3308_ MuI._3312_ MuI._3314_ vssd1 vssd1 vccd1 vccd1 MuI._3320_ sky130_fd_sc_hd__or3_1
X_10997_ _03736_ _03737_ _03553_ _03697_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__a211oi_1
XFILLER_15_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _05547_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__inv_2
XAuI._1074_ AuI._0199_ AuI._0200_ AuI._0284_ AuI._0223_ vssd1 vssd1 vccd1 vccd1 AuI._0285_
+ sky130_fd_sc_hd__a31o_1
XFILLER_204_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08664__A1 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4151_ MuI._3241_ MuI._3249_ vssd1 vssd1 vccd1 vccd1 MuI._3251_ sky130_fd_sc_hd__or2_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12667_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__nand2_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4082_ MuI._2858_ MuI._2859_ MuI._2863_ vssd1 vssd1 vccd1 vccd1 MuI._3182_ sky130_fd_sc_hd__a21o_1
XFILLER_175_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _04406_ _04407_ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or3_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _05460_ _05461_ _05439_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07120__A _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11549_ _02570_ _02741_ _04334_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and3b_1
XANTENNA__12961__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0927_ net29 AuI._0138_ vssd1 vssd1 vccd1 vccd1 AuI._0139_ sky130_fd_sc_hd__xnor2_4
XFILLER_100_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4984_ MuI._0723_ MuI._0716_ MuI._0722_ vssd1 vssd1 vccd1 vccd1 MuI._0726_ sky130_fd_sc_hd__and3_1
X_13219_ _06035_ _06046_ _06126_ _06043_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10481__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._0858_ net38 vssd1 vssd1 vccd1 vccd1 AuI._0078_ sky130_fd_sc_hd__inv_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6723_ MuI._2466_ MuI._2386_ MuI._2398_ vssd1 vssd1 vccd1 vccd1 MuI._2639_ sky130_fd_sc_hd__and3_1
XMuI._3935_ MuI._3033_ MuI._3034_ vssd1 vssd1 vccd1 vccd1 MuI._3035_ sky130_fd_sc_hd__and2b_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3866_ MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 MuI._2966_ sky130_fd_sc_hd__clkbuf_4
XMuI._6654_ MuI._1826_ MuI._2562_ vssd1 vssd1 vccd1 vccd1 MuI._2563_ sky130_fd_sc_hd__xor2_4
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08760_ _01374_ _01377_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._5605_ MuI._1370_ MuI._1374_ MuI._1376_ MuI._1400_ vssd1 vssd1 vccd1 vccd1 MuI._1409_
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07711_ _00318_ _00103_ _00327_ vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__or3_1
XFILLER_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3797_ MuI._2883_ MuI._2887_ MuI._2891_ MuI._2893_ MuI._2896_ vssd1 vssd1 vccd1
+ vccd1 MuI._2897_ sky130_fd_sc_hd__o221a_1
XMuI._6585_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2487_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08691_ _01066_ _01067_ _01117_ _01118_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__a22oi_2
XFILLER_93_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5536_ MuI._1327_ MuI._1328_ MuI._1323_ MuI._1326_ vssd1 vssd1 vccd1 vccd1 MuI._1333_
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07642_ _00257_ _00258_ _03163_ _00259_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__and4bb_1
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._416_ AuI.pe.significand\[21\] AuI.pe.significand\[23\] AuI.pe.significand\[22\]
+ AuI.pe.significand\[24\] vssd1 vssd1 vccd1 vccd1 AuI.pe._383_ sky130_fd_sc_hd__nor4b_1
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5467_ MuI._1250_ MuI._1251_ MuI._1256_ vssd1 vssd1 vccd1 vccd1 MuI._1257_ sky130_fd_sc_hd__a21o_1
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07573_ _06585_ _06583_ _06518_ _06562_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__and4_1
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4418_ MuI._2939_ MuI._2811_ MuI._3363_ MuI._0101_ vssd1 vssd1 vccd1 vccd1 MuI._0103_
+ sky130_fd_sc_hd__and4_1
XANTENNA_AuI.pe._683__A2 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ _01819_ _01818_ _01817_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10359__C _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5398_ MuI._1062_ MuI._1180_ vssd1 vssd1 vccd1 vccd1 MuI._1181_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4349_ MuI._1494_ MuI._2967_ vssd1 vssd1 vccd1 vccd1 MuI._0028_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI.pe._422__A AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _01859_ _01858_ _01640_ _01638_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o211a_1
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _01739_ _01738_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__and2b_1
XANTENNA_AuI._1285__B AuI._0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13400__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6019_ MuI._0878_ MuI._2797_ vssd1 vssd1 vccd1 vccd1 MuI._1864_ sky130_fd_sc_hd__nand2_1
XFILLER_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07030__A net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _00733_ _00742_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _00509_ _00510_ _00512_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__or3_1
XFILLER_116_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07007_ _05498_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11487__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10391__A _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__A2 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4305__A1 MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _01568_ _01569_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a21o_1
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07909_ _00524_ _00525_ _00526_ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__nand3_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _01495_ _01496_ _01505_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__and3_1
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ _03511_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__xnor2_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _03579_ _03580_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nand3_1
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10782_ _03504_ _03505_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand2_1
XFILLER_25_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12521_ _02849_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__inv_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _05303_ _05304_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__or2_1
XFILLER_185_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._831__C1 AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11403_ _04175_ _04177_ _02926_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XANTENNA__09071__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _05120_ _05122_ _05230_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o211ai_4
XFILLER_181_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09071__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11334_ _04101_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__xor2_4
XFILLER_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _03934_ _03936_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nand2_1
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11705__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ _03798_ _05456_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nand2_1
X_10216_ _02877_ _02898_ _02798_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21o_1
XFILLER_122_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11196_ _03951_ _03952_ _03948_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21o_1
XMuI._3720_ MuI._2814_ MuI._1142_ MuI._2786_ MuI._2352_ vssd1 vssd1 vccd1 vccd1 MuI._2820_
+ sky130_fd_sc_hd__and4_1
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09123__A2_N _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ _02823_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or2_1
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4847__A2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3504__C1 MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3651_ MuI._1791_ vssd1 vssd1 vccd1 vccd1 MuI._2517_ sky130_fd_sc_hd__buf_2
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10078_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__clkbuf_4
XMuI._6370_ MuI._2245_ MuI._2246_ MuI._2249_ vssd1 vssd1 vccd1 vccd1 MuI._2250_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3582_ MuI._1681_ MuI._1703_ vssd1 vssd1 vccd1 vccd1 MuI._1758_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13117__A _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5321_ MuI._1093_ MuI._1094_ MuI._1095_ vssd1 vssd1 vccd1 vccd1 MuI._1096_ sky130_fd_sc_hd__o21bai_1
XFILLER_75_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5252_ MuI.a_operand\[9\] MuI._3190_ MuI._2341_ MuI._3189_ vssd1 vssd1 vccd1
+ vccd1 MuI._1020_ sky130_fd_sc_hd__a22o_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1126_ AuI._0268_ AuI._0271_ AuI._0273_ AuI._0290_ AuI._0206_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0335_ sky130_fd_sc_hd__mux4_1
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4203_ MuI._3296_ MuI._3301_ MuI._3181_ vssd1 vssd1 vccd1 vccd1 MuI._3303_ sky130_fd_sc_hd__a21o_1
XANTENNA__06954__A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5183_ MuI._0940_ MuI._0943_ vssd1 vssd1 vccd1 vccd1 MuI._0945_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._3994__A MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ _02752_ _05489_ _05490_ _05592_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__a31o_4
XAuI._1057_ AuI._0266_ AuI._0267_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0268_ sky130_fd_sc_hd__mux2_1
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4134_ MuI._3232_ MuI._3222_ MuI._3229_ vssd1 vssd1 vccd1 vccd1 MuI._3234_ sky130_fd_sc_hd__and3_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07488__C _00105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__A1 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4065_ MuI._3161_ MuI._3163_ MuI._3164_ vssd1 vssd1 vccd1 vccd1 MuI._3165_ sky130_fd_sc_hd__or3_2
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12197__B2 AuI.result\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4783__B2 MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__A1 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _02032_ _02033_ _02024_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__o21ba_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4967_ MuI._0700_ MuI._0705_ MuI._0693_ MuI._0706_ vssd1 vssd1 vccd1 vccd1 MuI._0707_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09861_ _02479_ _02492_ _02516_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__and3_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6706_ MuI._2615_ MuI._2619_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2620_ sky130_fd_sc_hd__mux2_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08112__C _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3918_ MuI._2938_ MuI._3012_ MuI._3017_ vssd1 vssd1 vccd1 vccd1 MuI._3018_ sky130_fd_sc_hd__o21ai_1
X_08812_ _01391_ _01392_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4898_ MuI._0436_ MuI._0630_ vssd1 vssd1 vccd1 vccd1 MuI._0631_ sky130_fd_sc_hd__nand2_1
X_09792_ _02393_ _02403_ _02406_ _02441_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__or4bb_1
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6637_ MuI._1760_ MuI._2543_ vssd1 vssd1 vccd1 vccd1 MuI._2544_ sky130_fd_sc_hd__xnor2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3849_ MuI._2945_ MuI._2948_ vssd1 vssd1 vccd1 vccd1 MuI._2949_ sky130_fd_sc_hd__and2_1
X_08743_ _01359_ _01360_ _06608_ _00301_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__and4bb_1
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6568_ MuI._2426_ MuI._2443_ vssd1 vssd1 vccd1 vccd1 MuI._2468_ sky130_fd_sc_hd__nand2_1
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__D _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08674_ _01278_ _01290_ _01289_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__a21o_1
XFILLER_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07670__D _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5519_ MuI._2967_ MuI._0245_ MuI._1300_ MuI._1299_ vssd1 vssd1 vccd1 vccd1 MuI._1314_
+ sky130_fd_sc_hd__a31o_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07025__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07625_ _00240_ _00241_ _00242_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__and3_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6499_ MuI._2378_ MuI._2391_ MuI._2379_ vssd1 vssd1 vccd1 vccd1 MuI._2392_ sky130_fd_sc_hd__o21bai_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__D _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5263__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07556_ _06651_ _06653_ _06652_ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12424__A2 _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06864__A _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10435__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6212__A1 MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10386__A _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07487_ _00103_ _00104_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__or2_2
XFILLER_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _01765_ _01768_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__and3_1
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09157_ _01772_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__or2b_1
XFILLER_175_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08108_ _00722_ _00723_ _00724_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _01701_ _01705_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _00255_ _00256_ _00368_ _00369_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__a22oi_2
XFILLER_135_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09356__A2 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _03780_ _03794_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nand3_2
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10001_ _02650_ _02654_ _02653_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _02862_ _05906_ _05981_ _02808_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__a22o_1
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6174__B MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0915__A0 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _03596_ _03597_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__o211a_1
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _04675_ _04676_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a21o_1
XFILLER_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ _00058_ _00002_ _03560_ _03562_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__nand4_1
XANTENNA__06774__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0822__B net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _02767_ _03302_ _02498_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A2 _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12504_ _04994_ _02728_ _02732_ AuI.result\[16\] vssd1 vssd1 vccd1 vccd1 _05362_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_AuI._0861__A2_N net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13484_ _02744_ _02812_ _02945_ _05917_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a221o_1
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _03379_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xor2_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12179__B2 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12435_ _05269_ _05286_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__nand2_1
XFILLER_154_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__and2_1
XFILLER_181_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5714__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5870_ MuI._1682_ MuI._1683_ MuI._1698_ MuI._1699_ vssd1 vssd1 vccd1 vccd1 MuI._1700_
+ sky130_fd_sc_hd__or4_1
X_11317_ _04074_ _04084_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xor2_1
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _02752_ _05019_ _05020_ _05139_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__a31o_2
XAuI.pe._750_ AuI.pe._024_ AuI.pe._293_ vssd1 vssd1 vccd1 vccd1 AuI.pe._294_ sky130_fd_sc_hd__or2_1
XMuI._4821_ MuI._0502_ MuI._0544_ MuI._0545_ vssd1 vssd1 vccd1 vccd1 MuI._0546_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output75_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._583__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _02707_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1675_ net29 AuI._0126_ AuI._0699_ AuI._0024_ vssd1 vssd1 vccd1 vccd1 AuI.result\[31\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07697__A_N _00313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._681_ AuI.pe._071_ AuI.pe._150_ AuI.pe._173_ AuI.pe.significand\[4\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._229_ sky130_fd_sc_hd__a22o_1
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4752_ MuI._0457_ MuI._0462_ MuI._0464_ vssd1 vssd1 vccd1 vccd1 MuI._0470_ sky130_fd_sc_hd__or3_1
XFILLER_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11179_ _03926_ _03934_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__nand3_1
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3703_ MuI._2638_ vssd1 vssd1 vccd1 vccd1 MuI._2803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4683_ MuI._0385_ MuI._0389_ MuI._0391_ vssd1 vssd1 vccd1 vccd1 MuI._0395_ sky130_fd_sc_hd__o21ai_1
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3634_ MuI._2319_ vssd1 vssd1 vccd1 vccd1 MuI._2330_ sky130_fd_sc_hd__buf_2
XMuI._6422_ MuI._2241_ MuI._2306_ vssd1 vssd1 vccd1 vccd1 MuI._2307_ sky130_fd_sc_hd__or2_1
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08586__D _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08858__A1 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08858__B2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6353_ MuI._2207_ MuI._2230_ vssd1 vssd1 vccd1 vccd1 MuI._2232_ sky130_fd_sc_hd__nor2_1
XMuI._3565_ MuI._1230_ MuI._1560_ vssd1 vssd1 vccd1 vccd1 MuI._1571_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10665__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10665__B2 _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5304_ MuI._2898_ MuI._0112_ MuI._1075_ MuI._1077_ vssd1 vssd1 vccd1 vccd1 MuI._1078_
+ sky130_fd_sc_hd__a31oi_2
XMuI._6284_ MuI._2140_ MuI._2141_ vssd1 vssd1 vccd1 vccd1 MuI._2156_ sky130_fd_sc_hd__and2b_1
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07410_ net120 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__clkbuf_4
XMuI._3496_ MuI._0801_ MuI._0471_ vssd1 vssd1 vccd1 vccd1 MuI._0812_ sky130_fd_sc_hd__nand2_1
XANTENNA__12406__A2 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ _01004_ _01006_ _01005_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a21o_1
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5235_ MuI._1000_ MuI._1001_ vssd1 vssd1 vccd1 vccd1 MuI._1002_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _06556_ _06557_ _06573_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__nand3_1
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1109_ AuI._0261_ AuI._0309_ AuI._0318_ vssd1 vssd1 vccd1 vccd1 AuI._0319_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._5709__A MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08086__A2 _00702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._1331__A0 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5166_ MuI._0905_ MuI._0924_ MuI._0925_ vssd1 vssd1 vccd1 vccd1 MuI._0926_ sky130_fd_sc_hd__and3_1
XFILLER_149_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07272_ _06558_ _06572_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__xor2_1
XFILLER_192_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3874__D MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4117_ MuI._2919_ MuI._2528_ MuI._2539_ MuI._2800_ vssd1 vssd1 vccd1 vccd1 MuI._3217_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_177_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _01291_ _01292_ _01294_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a21oi_2
XMuI._5097_ MuI._0477_ MuI._3402_ MuI._3396_ MuI._0327_ vssd1 vssd1 vccd1 vccd1 MuI._0850_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_192_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4048_ MuI._3056_ MuI._3126_ MuI._3145_ MuI._3146_ vssd1 vssd1 vccd1 vccd1 MuI._3148_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07597__A1 _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__A2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07597__B2 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6259__B MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5181__A1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09913_ _02551_ _02571_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5181__B2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5999_ MuI._3037_ MuI._3156_ vssd1 vssd1 vccd1 vccd1 MuI._1842_ sky130_fd_sc_hd__and2_1
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1398__B1 AuI._0586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _02462_ _02461_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__and2b_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06859__A _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09775_ _02407_ _02408_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__nand3_2
X_06987_ _05284_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[20\] sky130_fd_sc_hd__clkbuf_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _06519_ _06515_ net6 net7 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and4_1
XFILLER_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12645__A2 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _01214_ _01274_ _01272_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a21o_1
XFILLER_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07608_ _00223_ _00224_ _00214_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__a21o_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08588_ _00462_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__buf_4
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _00151_ _00154_ _00152_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13204__B _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1322__A0 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11081__A1 _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07285__B1 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _00164_ _06500_ _03082_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__and3_1
XFILLER_167_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4242__B MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _01812_ _01824_ _01823_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a21o_1
XFILLER_182_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _02905_ _02959_ _00423_ _05198_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__nand4_1
XANTENNA__10844__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _05052_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12030__B1 _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12581__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _04979_ _04980_ _04849_ _04941_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__o211ai_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ _02879_ _02886_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__and2_1
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _00216_ _05820_ _03444_ _00217_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a22oi_1
XFILLER_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09734__C1 _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11033_ _03612_ _03614_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__nand2_1
XFILLER_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1460_ AuI._0376_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0646_ sky130_fd_sc_hd__and2_1
XFILLER_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07872__B _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12884__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06769__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0817__B net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__B _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1391_ AuI._0581_ AuI._0573_ AuI._0567_ vssd1 vssd1 vccd1 vccd1 AuI._0582_ sky130_fd_sc_hd__a21o_1
XFILLER_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6185__A MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3486__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12984_ _03497_ _05713_ _05790_ _05789_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__a31o_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ _04554_ _04598_ _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__o211a_2
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0833__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._504__B AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _04672_ _04673_ _04674_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a21o_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10817_ _03360_ _03362_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__nand2_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5020_ MuI._0760_ MuI._0763_ MuI._0764_ MuI._0611_ vssd1 vssd1 vccd1 vccd1 MuI._0765_
+ sky130_fd_sc_hd__o211a_1
X_11797_ _04469_ _04471_ _04600_ _04601_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a211o_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10748_ _03272_ _03274_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11252__A1_N _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ _06376_ _06379_ _06380_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__or4_1
X_10679_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nor2_1
XFILLER_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12418_ _05154_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__xnor2_1
XFILLER_154_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13398_ FuI.Integer\[28\] _06056_ _02745_ _06016_ _06311_ vssd1 vssd1 vccd1 vccd1
+ _06312_ sky130_fd_sc_hd__a221o_1
XANTENNA__08224__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07766__C net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5922_ MuI._1649_ MuI._1708_ MuI._1707_ vssd1 vssd1 vccd1 vccd1 MuI._1757_ sky130_fd_sc_hd__a21boi_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _05193_ _05191_ _05192_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nand3_2
XFILLER_141_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._802_ AuI.pe._330_ AuI.pe._341_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[2\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5853_ MuI._1581_ MuI._1668_ MuI._1679_ MuI._1680_ vssd1 vssd1 vccd1 vccd1 MuI._1682_
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._556__A1 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._733_ AuI.pe._102_ AuI.pe._164_ AuI.pe._397_ AuI.pe._072_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._278_ sky130_fd_sc_hd__a22o_1
XMuI._4804_ MuI._0491_ MuI._0524_ MuI._0525_ MuI._0527_ vssd1 vssd1 vccd1 vccd1 MuI._0528_
+ sky130_fd_sc_hd__and4_1
X_06910_ _04456_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__clkbuf_4
XMuI._5784_ MuI._1508_ MuI._1510_ vssd1 vssd1 vccd1 vccd1 MuI._1606_ sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1658_ AuI._0604_ AuI._0710_ vssd1 vssd1 vccd1 vccd1 AuI._0012_ sky130_fd_sc_hd__nand2_1
X_07890_ net112 _03593_ _06431_ _00287_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__and4_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._664_ AuI.pe.significand\[7\] AuI.pe._197_ AuI.pe._071_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._213_ sky130_fd_sc_hd__and3b_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4735_ MuI._0321_ MuI._0316_ vssd1 vssd1 vccd1 vccd1 MuI._0452_ sky130_fd_sc_hd__and2_1
XANTENNA__08597__C _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06841_ net60 vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__buf_2
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1589_ AuI._0761_ AuI._0762_ vssd1 vssd1 vccd1 vccd1 AuI._0763_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11735__D _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._595_ AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 AuI.pe._149_ sky130_fd_sc_hd__inv_2
XMuI._4666_ MuI.a_operand\[20\] MuI.a_operand\[19\] MuI.b_operand\[1\] MuI.b_operand\[0\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0376_ sky130_fd_sc_hd__and4_1
X_09560_ _02377_ _00301_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__nand2_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06772_ _02970_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and3_1
XFILLER_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6405_ MuI._2285_ MuI._2278_ MuI._2288_ vssd1 vssd1 vccd1 vccd1 MuI._2289_ sky130_fd_sc_hd__a21o_1
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3617_ MuI._1780_ MuI._2132_ vssd1 vssd1 vccd1 vccd1 MuI._2143_ sky130_fd_sc_hd__and2b_1
X_08511_ _01060_ _01062_ _01127_ _01128_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a211oi_4
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4597_ MuI._0220_ MuI._0222_ vssd1 vssd1 vccd1 vccd1 MuI._0300_ sky130_fd_sc_hd__xnor2_1
X_09491_ _02110_ _02111_ _02116_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__nand3_1
XFILLER_24_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6336_ MuI._2211_ MuI._2212_ vssd1 vssd1 vccd1 vccd1 MuI._2213_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3548_ MuI._0889_ MuI._0801_ vssd1 vssd1 vccd1 vccd1 MuI._1384_ sky130_fd_sc_hd__nand2_1
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _01057_ _01058_ _01059_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a21o_1
XFILLER_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6267_ MuI._2135_ MuI._2136_ vssd1 vssd1 vccd1 vccd1 MuI._2137_ sky130_fd_sc_hd__nor2_1
XMuI._3479_ MuI._0614_ vssd1 vssd1 vccd1 vccd1 MuI._0625_ sky130_fd_sc_hd__clkbuf_4
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07303__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__A2 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _00988_ _00989_ _00990_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__or3_1
XFILLER_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5218_ MuI._0975_ MuI._0981_ MuI._0952_ MuI._0953_ vssd1 vssd1 vccd1 vccd1 MuI._0983_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08118__B _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07324_ _06583_ _06623_ _05187_ _06585_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__a22o_1
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6198_ MuI._2059_ MuI._2060_ vssd1 vssd1 vccd1 vccd1 MuI._2061_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07806__A2 _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4062__B MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5149_ MuI._2765_ MuI._2885_ MuI._2881_ MuI._2484_ vssd1 vssd1 vccd1 vccd1 MuI._0907_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ _06553_ _06554_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nand3_2
XFILLER_118_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07186_ _06470_ _06468_ _06467_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o21ai_1
XFILLER_133_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08134__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B1 _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__B2 _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12315__A1 _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11495__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__B2 _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07692__B net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _02436_ _02437_ _02429_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__o21ba_1
XFILLER_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5848__A1_N MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ _02404_ _02405_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__nor2_1
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._605__A AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _01200_ _01326_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__xor2_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11826__B1 _04623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _02014_ _02015_ _02016_ _01996_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ _04513_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__nand3_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4417__B1 MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07213__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5349__A MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ _00502_ _04607_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__nand2_1
XFILLER_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _02741_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__buf_4
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11582_ _04367_ _04368_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__or2_1
XFILLER_156_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13321_ _06227_ _06172_ _06230_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__nor3_1
XANTENNA_MuI._4403__D MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10533_ _03220_ _03238_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__and3_1
XAuI._0960_ net44 net12 AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0172_ sky130_fd_sc_hd__mux2_1
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09094__A1_N _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13252_ _06158_ _06159_ _04635_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__mux2_1
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10464_ _03162_ _03164_ _03159_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a21o_1
XFILLER_171_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0891_ AuI._0103_ AuI._0106_ AuI._0109_ AuI._0110_ vssd1 vssd1 vccd1 vccd1 AuI._0111_
+ sky130_fd_sc_hd__o31a_1
XFILLER_182_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12203_ _04906_ _04937_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__or2b_1
XANTENNA__08758__B1 _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _02645_ _06089_ _04159_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__a21oi_1
X_10395_ _00792_ _00793_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__and2b_1
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12134_ _00283_ _05198_ _04960_ _04962_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nand4_2
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1512_ AuI._0116_ AuI._0697_ vssd1 vssd1 vccd1 vccd1 AuI._0698_ sky130_fd_sc_hd__or2_1
X_12065_ _04161_ _04884_ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _03324_ _00445_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__nand2_1
XANTENNA__10868__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09722__A2 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1443_ AuI._0515_ AuI._0519_ AuI._0622_ AuI._0628_ vssd1 vssd1 vccd1 vccd1 AuI._0629_
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__10868__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4520_ MuI._0213_ MuI._0090_ MuI._0214_ vssd1 vssd1 vccd1 vccd1 MuI._0215_ sky130_fd_sc_hd__or3_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1374_ net17 net49 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0566_ sky130_fd_sc_hd__mux2_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4451_ MuI._0016_ MuI._0138_ vssd1 vssd1 vccd1 vccd1 MuI._0139_ sky130_fd_sc_hd__or2b_1
XFILLER_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__B1 _01350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _02801_ _05273_ _02806_ _02807_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__o31ai_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4382_ MuI._0042_ MuI._0045_ vssd1 vssd1 vccd1 vccd1 MuI._0064_ sky130_fd_sc_hd__or2b_1
XFILLER_61_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13125__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _04576_ _04578_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nand2_1
XANTENNA__11293__A1 _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12490__B1 _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _05603_ _05782_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o21a_1
XMuI._6121_ MuI._1970_ MuI._1975_ vssd1 vssd1 vccd1 vccd1 MuI._1976_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _05970_ _04655_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._4163__A MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6052_ MuI._3067_ MuI._1899_ vssd1 vssd1 vccd1 vccd1 MuI._1900_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07249__B1 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5003_ MuI._0555_ MuI._0744_ MuI._0745_ vssd1 vssd1 vccd1 vccd1 MuI._0747_ sky130_fd_sc_hd__nand3_1
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ _05853_ _02042_ _02151_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__and3_1
XFILLER_162_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08749__B1 _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12545__A1 _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12545__B2 _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5905_ MuI._0755_ MuI._0756_ vssd1 vssd1 vccd1 vccd1 MuI._1739_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07793__A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__B1 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _01470_ _01471_ _01480_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and3_1
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5836_ MuI._1660_ MuI._1662_ vssd1 vssd1 vccd1 vccd1 MuI._1663_ sky130_fd_sc_hd__xor2_1
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07942_ _00536_ _00543_ _00544_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__nand3_1
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._716_ AuI.pe.significand\[20\] AuI.pe.significand\[23\] AuI.pe._035_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._262_ sky130_fd_sc_hd__a21o_1
XANTENNA__12204__A _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08401__B _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5767_ MuI._1585_ MuI._1586_ vssd1 vssd1 vccd1 vccd1 MuI._1587_ sky130_fd_sc_hd__nor2_1
X_07873_ _00486_ _00489_ _00490_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__nand3_2
XAuI.pe._647_ AuI.pe._370_ AuI.pe._374_ vssd1 vssd1 vccd1 vccd1 AuI.pe._197_ sky130_fd_sc_hd__nor2_4
XFILLER_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4718_ MuI._0430_ MuI._0432_ vssd1 vssd1 vccd1 vccd1 MuI._0433_ sky130_fd_sc_hd__or2_1
XFILLER_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09612_ _02245_ _02246_ _02247_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a21bo_1
X_06824_ net112 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__buf_2
XMuI._5698_ MuI._1508_ MuI._1509_ MuI._1507_ vssd1 vssd1 vccd1 vccd1 MuI._1511_ sky130_fd_sc_hd__a21bo_1
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4057__B MuI._3156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._578_ AuI.pe._132_ vssd1 vssd1 vccd1 vccd1 AuI.pe._133_ sky130_fd_sc_hd__buf_2
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4649_ MuI._0354_ MuI._0356_ vssd1 vssd1 vccd1 vccd1 MuI._0357_ sky130_fd_sc_hd__or2b_1
X_09543_ _02528_ _04111_ _02055_ _02056_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XANTENNA__11762__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06755_ net41 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__buf_4
XANTENNA__10659__A _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09474_ _06494_ _06495_ _00084_ _04574_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3870__A1 MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06686_ _02042_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__buf_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6319_ MuI._2155_ MuI._2193_ vssd1 vssd1 vccd1 vccd1 MuI._2194_ sky130_fd_sc_hd__or2b_1
XANTENNA__07033__A _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08425_ _01038_ _01039_ _01042_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__nand3_1
XFILLER_197_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08356_ _06491_ _05241_ _05305_ _06492_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06872__A _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08790__C _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07307_ net121 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__buf_4
X_08287_ _00874_ _00902_ _00903_ _00904_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__nand4_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07238_ _06535_ _06536_ _06538_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or3_1
XFILLER_192_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._768__A1 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12536__A1 AuI.result\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__B _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07169_ _06469_ _02194_ net22 _05627_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__and4_1
XFILLER_106_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10180_ _02858_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__nand2_2
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5678__A2 MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12114__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09126__C _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11953__A _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12821_ _05698_ _05699_ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__o21a_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1090_ AuI._0139_ AuI._0298_ AuI._0299_ vssd1 vssd1 vccd1 vccd1 AuI._0301_ sky130_fd_sc_hd__o21bai_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _05624_ _05625_ _05535_ _05539_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o211ai_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12472__B1 _05308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ _04373_ _04378_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__nand2_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _05551_ _05552_ _05511_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__o21a_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _04365_ _04249_ _04424_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o211ai_4
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11565_ _04542_ _02728_ _02938_ AuI.result\[9\] vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09640__A1 _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09640__B2 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ _06211_ _06213_ _06214_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__or3_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _02840_ _06561_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._759__A1 AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0943_ net55 net23 AuI._0121_ vssd1 vssd1 vccd1 vccd1 AuI._0155_ sky130_fd_sc_hd__mux2_1
XANTENNA__07651__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ _04272_ _04276_ _04277_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__nand3_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13235_ _05595_ _02941_ _02837_ _03306_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__o22ai_1
XFILLER_6_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10447_ _03145_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10538__B1 _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0874_ net49 AuI._0027_ AuI._0033_ vssd1 vssd1 vccd1 vccd1 AuI._0094_ sky130_fd_sc_hd__a21oi_1
XMuI._3951_ MuI._3049_ MuI._3050_ vssd1 vssd1 vccd1 vccd1 MuI._3051_ sky130_fd_sc_hd__and2b_1
XFILLER_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11847__B _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _06063_ _06071_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__nand2_1
XANTENNA__10936__A1_N _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ _06560_ _03071_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._6638__A MuI._1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6670_ MuI._2574_ MuI._2579_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2580_ sky130_fd_sc_hd__mux2_1
X_12117_ _06439_ _00197_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__nand2_1
XMuI._3882_ MuI._2978_ MuI._2979_ MuI._2980_ vssd1 vssd1 vccd1 vccd1 MuI._2982_ sky130_fd_sc_hd__a21o_1
XFILLER_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13097_ _02643_ _02638_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__or2b_1
XFILLER_123_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5621_ MuI._1421_ MuI._1423_ MuI._1425_ vssd1 vssd1 vccd1 vccd1 MuI._1426_ sky130_fd_sc_hd__o21a_1
XANTENNA__07118__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ _04870_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__xnor2_1
XAuI.pe._501_ AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 AuI.pe._062_ sky130_fd_sc_hd__buf_2
XMuI._5552_ MuI._3268_ MuI._0445_ vssd1 vssd1 vccd1 vccd1 MuI._1350_ sky130_fd_sc_hd__nand2_1
XAuI._1426_ AuI._0253_ AuI._0611_ vssd1 vssd1 vccd1 vccd1 AuI._0612_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._432_ AuI.pe._367_ AuI.pe._384_ AuI.pe._387_ vssd1 vssd1 vccd1 vccd1 AuI.pe._399_
+ sky130_fd_sc_hd__and3_2
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06957__A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4503_ MuI._0172_ MuI._0178_ vssd1 vssd1 vccd1 vccd1 MuI._0197_ sky130_fd_sc_hd__or2b_1
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5483_ MuI._1265_ MuI._1266_ vssd1 vssd1 vccd1 vccd1 MuI._1275_ sky130_fd_sc_hd__and2_1
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__B _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1357_ AuI._0549_ AuI._0550_ vssd1 vssd1 vccd1 vccd1 AuI._0551_ sky130_fd_sc_hd__xor2_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4434_ MuI._0064_ MuI._0066_ MuI._0068_ vssd1 vssd1 vccd1 vccd1 MuI._0121_ sky130_fd_sc_hd__a21o_1
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11266__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__B2 _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1288_ AuI._0212_ AuI._0261_ vssd1 vssd1 vccd1 vccd1 AuI._0487_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4605__B MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4365_ MuI._0042_ MuI._0045_ vssd1 vssd1 vccd1 vccd1 MuI._0046_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12694__A _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6104_ MuI._1926_ MuI._1957_ vssd1 vssd1 vccd1 vccd1 MuI._1958_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08210_ _06463_ net19 _05434_ _02107_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__a22oi_2
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4296_ MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 MuI._3396_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11018__A1 _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ _01743_ _01745_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__nand2_1
XANTENNA__11018__B2 _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06692__A _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6035_ MuI._3103_ MuI._3119_ vssd1 vssd1 vccd1 vccd1 MuI._1882_ sky130_fd_sc_hd__or2b_1
XFILLER_193_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08141_ _00756_ _00757_ _00758_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__or3_1
XFILLER_174_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08072_ _00502_ _03993_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__nand2_1
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12518__A1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _05671_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and3_1
XFILLER_162_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout107_A net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08412__A _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6868_ MuI._2735_ MuI._2769_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[26\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08974_ _01457_ _01459_ _01458_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nand3_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5819_ MuI._1642_ MuI._1643_ vssd1 vssd1 vccd1 vccd1 MuI._1644_ sky130_fd_sc_hd__and2b_1
XANTENNA__07028__A _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _00540_ _00542_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__or2b_1
XMuI._6799_ MuI._2719_ MuI._2720_ MuI._2721_ vssd1 vssd1 vccd1 vccd1 MuI._2722_ sky130_fd_sc_hd__a21bo_1
XFILLER_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__A _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ _00204_ _00207_ _00472_ _00473_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a211oi_1
XANTENNA__06867__A _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06807_ _03346_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__and3_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4218__D MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _00394_ _00404_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__xor2_1
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3700__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ _02068_ _02072_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a21bo_1
X_06738_ _02042_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__clkbuf_2
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4515__B MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _02066_ _02076_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__or3_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08408_ _02723_ _04660_ _01024_ _01025_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__a31o_1
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08009__D _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _01917_ _01916_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__and2b_1
XANTENNA__10480__A2 _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._112_ FuI._023_ FuI._054_ vssd1 vssd1 vccd1 vccd1 FuI._024_ sky130_fd_sc_hd__nor2_1
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08339_ _00829_ _00827_ _00828_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__or3_1
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10768__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _02987_ _06613_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__nand4_1
XANTENNA_MuI._5346__B MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__A1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10301_ _00695_ _00697_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nand2_1
XFILLER_125_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _03916_ _04043_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__nand3_2
X_13020_ _05864_ _05832_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a21o_1
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4571__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10232_ _03755_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__inv_2
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5362__A MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _02830_ _02833_ _02837_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5520__A1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5520__B2 MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input37_A b_operand[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10094_ _02302_ _04122_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13485__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08976__B _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06777__A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08361__A1 _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09153__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08361__B2 _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1211_ AuI._0412_ AuI._0414_ AuI._0415_ vssd1 vssd1 vccd1 vccd1 AuI._0416_ sky130_fd_sc_hd__and3_1
XFILLER_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4087__A1 MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4706__A MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3610__A MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0960__A1 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1142_ AuI._0177_ AuI._0183_ AuI._0310_ AuI._0311_ AuI._0274_ AuI._0276_ vssd1
+ vssd1 vccd1 vccd1 AuI._0350_ sky130_fd_sc_hd__mux4_1
X_12804_ _05684_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996_ _03553_ _03697_ _03736_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__o211a_1
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12735_ _05608_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__xnor2_1
XAuI._1073_ net63 net62 net31 net30 AuI._0174_ AuI._0124_ vssd1 vssd1 vccd1 vccd1
+ AuI._0284_ sky130_fd_sc_hd__mux4_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08664__A2 _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4150_ MuI._3241_ MuI._3249_ vssd1 vssd1 vccd1 vccd1 MuI._3250_ sky130_fd_sc_hd__nand2_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__A_N _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12666_ _05533_ _05534_ _05529_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__a21o_1
XFILLER_129_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3598__B1 MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4081_ MuI._2960_ MuI._3180_ vssd1 vssd1 vccd1 vccd1 MuI._3181_ sky130_fd_sc_hd__xor2_1
X_11617_ _00088_ _03047_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__nand2_1
X_12597_ _05439_ _05460_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XFILLER_168_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11548_ _02546_ _02569_ _04157_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__a21bo_1
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12961__B _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11858__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0926_ AuI.AddBar_Sub net61 vssd1 vssd1 vccd1 vccd1 AuI._0138_ sky130_fd_sc_hd__xor2_4
X_11479_ _04257_ _04258_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__xor2_2
XANTENNA__13173__A1 _04211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ _06041_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__clkinv_2
XMuI._4983_ MuI._0716_ MuI._0722_ MuI._0723_ vssd1 vssd1 vccd1 vccd1 MuI._0725_ sky130_fd_sc_hd__a21oi_4
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0857_ AuI._0069_ AuI._0072_ AuI._0073_ AuI._0076_ vssd1 vssd1 vccd1 vccd1 AuI._0077_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_140_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10481__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6722_ MuI._2386_ MuI._2398_ MuI._2466_ vssd1 vssd1 vccd1 vccd1 MuI._2637_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3934_ MuI._3027_ MuI._3031_ MuI._3032_ vssd1 vssd1 vccd1 vccd1 MuI._3034_ sky130_fd_sc_hd__or3b_1
XFILLER_152_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__or2_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6653_ MuI._1827_ MuI._1828_ MuI._2560_ vssd1 vssd1 vccd1 vccd1 MuI._2562_ sky130_fd_sc_hd__o21a_1
XFILLER_100_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3865_ MuI._2962_ MuI._2963_ MuI._2961_ vssd1 vssd1 vccd1 vccd1 MuI._2965_ sky130_fd_sc_hd__a21bo_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._5604_ MuI._1402_ MuI._1405_ MuI._1407_ vssd1 vssd1 vccd1 vccd1 MuI._1408_ sky130_fd_sc_hd__nand3_1
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _00318_ _00103_ _00327_ vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__o21ai_2
XFILLER_211_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6584_ MuI._2485_ vssd1 vssd1 vccd1 vccd1 MuI._2486_ sky130_fd_sc_hd__clkbuf_4
XMuI._3796_ MuI._2894_ MuI._2895_ vssd1 vssd1 vccd1 vccd1 MuI._2896_ sky130_fd_sc_hd__and2_1
X_08690_ _01304_ _01305_ _01306_ _01307_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__nand4_1
XANTENNA__06687__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5535_ MuI._1287_ MuI._1291_ MuI._1294_ MuI._1330_ vssd1 vssd1 vccd1 vccd1 MuI._1332_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09063__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1409_ AuI._0410_ AuI._0498_ vssd1 vssd1 vccd1 vccd1 AuI._0598_ sky130_fd_sc_hd__or2_2
X_07641_ _00074_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__buf_4
XAuI.pe._415_ AuI.pe.significand\[16\] vssd1 vssd1 vccd1 vccd1 AuI.pe._382_ sky130_fd_sc_hd__inv_2
XANTENNA_MuI._4616__A MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5466_ MuI._1253_ MuI._1254_ MuI._1255_ vssd1 vssd1 vccd1 vccd1 MuI._1256_ sky130_fd_sc_hd__o21bai_1
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _02658_ _05252_ _05316_ _02593_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__a22oi_2
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4417_ MuI._2813_ MuI._3363_ MuI._0101_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._0102_
+ sky130_fd_sc_hd__a22oi_1
X_09311_ _01819_ _01817_ _01818_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__or3_1
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5397_ MuI._1172_ MuI._1178_ MuI._1179_ vssd1 vssd1 vccd1 vccd1 MuI._1180_ sky130_fd_sc_hd__o21a_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10359__D _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4348_ MuI._0024_ MuI._0026_ vssd1 vssd1 vccd1 vccd1 MuI._0027_ sky130_fd_sc_hd__or2_1
X_09242_ _01638_ _01640_ _01858_ _01859_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a211oi_2
XFILLER_61_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4888__A1_N MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07311__A _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4279_ MuI._3357_ MuI._3378_ vssd1 vssd1 vccd1 vccd1 MuI._3379_ sky130_fd_sc_hd__or2_1
X_09173_ _02851_ _04046_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4351__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6018_ MuI._0878_ MuI._2789_ MuI._3107_ vssd1 vssd1 vccd1 vccd1 MuI._1863_ sky130_fd_sc_hd__and3_1
X_08124_ _00740_ _00741_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__or2b_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _00441_ _00475_ _00474_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__o21bai_2
XFILLER_174_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ net21 vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11487__B _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10391__B _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5613__C MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _01570_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07908_ _00523_ _00522_ _00370_ _00255_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__o211ai_4
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _01495_ _01496_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a21oi_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09540__B1 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07839_ _03271_ _04509_ _00035_ _03217_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__a22o_1
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _03152_ _06580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__and2_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _02127_ _02128_ _02135_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10781_ _03504_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__or2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12520_ _02752_ _05264_ _05265_ _05378_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__a31o_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net61 _05058_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4261__A MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _02879_ _02886_ _02757_ _02887_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__a31o_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ _05228_ _05229_ _05114_ _05145_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__a211o_1
XFILLER_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09071__A2 _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ _02965_ _04596_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nand2_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _03945_ _03946_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__or4_2
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11166__B1 _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__A2 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _05894_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__nor2_1
XFILLER_79_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10215_ _02897_ _02795_ _02793_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__o21bai_1
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11195_ _03948_ _03951_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__nand3_1
XFILLER_122_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _03680_ _05853_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__and2b_1
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3650_ MuI._2473_ MuI._2495_ vssd1 vssd1 vccd1 vccd1 MuI._2506_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4139__C MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10077_ _02020_ _06023_ _02075_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__and3_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3581_ MuI._1648_ MuI._1714_ MuI._1736_ vssd1 vssd1 vccd1 vccd1 MuI._1747_ sky130_fd_sc_hd__a21oi_1
XFILLER_208_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5320_ MuI._2785_ MuI._2341_ MuI._3262_ MuI._0020_ vssd1 vssd1 vccd1 vccd1 MuI._1095_
+ sky130_fd_sc_hd__and4_1
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11543__A1_N _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5251_ MuI._2873_ MuI._2785_ MuI._2875_ MuI._3349_ vssd1 vssd1 vccd1 vccd1 MuI._1019_
+ sky130_fd_sc_hd__nand4_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09611__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1125_ AuI._0263_ AuI._0333_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0334_ sky130_fd_sc_hd__o21a_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979_ _03486_ _00059_ _03717_ _03718_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a22o_1
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13091__B1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4202_ MuI._3181_ MuI._3296_ MuI._3301_ vssd1 vssd1 vccd1 vccd1 MuI._3302_ sky130_fd_sc_hd__and3_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5182_ MuI._0941_ MuI._0942_ vssd1 vssd1 vccd1 vccd1 MuI._0943_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._3994__B MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _05570_ _05571_ _05577_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__a211o_1
XANTENNA__07845__B1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A1 _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1056_ AuI._0164_ AuI._0169_ AuI._0216_ vssd1 vssd1 vccd1 vccd1 AuI._0267_ sky130_fd_sc_hd__and3_1
XFILLER_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4133_ MuI._3222_ MuI._3229_ MuI._3232_ vssd1 vssd1 vccd1 vccd1 MuI._3233_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07131__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12649_ _05515_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__xnor2_1
XMuI._4064_ MuI._2905_ MuI._2904_ MuI._2879_ vssd1 vssd1 vccd1 vccd1 MuI._3164_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13394__A1 _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4783__A2 MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__B2 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06970__A _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0909_ AuI._0111_ AuI._0114_ AuI._0117_ AuI._0118_ vssd1 vssd1 vccd1 vccd1 AuI._0128_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6098__A MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3515__A MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4966_ MuI._0682_ MuI._0689_ MuI._0692_ vssd1 vssd1 vccd1 vccd1 MuI._0706_ sky130_fd_sc_hd__nand3_1
X_09860_ _02511_ _02513_ _02515_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a21oi_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6705_ MuI._2366_ MuI._2618_ vssd1 vssd1 vccd1 vccd1 MuI._2619_ sky130_fd_sc_hd__xor2_2
XFILLER_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3917_ MuI._3015_ MuI._3016_ vssd1 vssd1 vccd1 vccd1 MuI._3017_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _01427_ _01428_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__nand2_1
XANTENNA__08112__D _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4897_ MuI._0433_ MuI._0435_ vssd1 vssd1 vccd1 vccd1 MuI._0630_ sky130_fd_sc_hd__or2_1
X_09791_ _02436_ _02438_ _02439_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__o211a_1
XFILLER_98_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6636_ MuI._1712_ MuI._2537_ MuI._1762_ vssd1 vssd1 vccd1 vccd1 MuI._2543_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3848_ MuI._2946_ MuI._2947_ vssd1 vssd1 vccd1 vccd1 MuI._2948_ sky130_fd_sc_hd__xor2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _02797_ _00074_ _00090_ _02754_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__a22oi_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6567_ MuI._2386_ MuI._2398_ MuI._2460_ MuI._2466_ vssd1 vssd1 vccd1 vccd1 MuI._2467_
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3779_ MuI._2870_ MuI._2878_ vssd1 vssd1 vccd1 vccd1 MuI._2879_ sky130_fd_sc_hd__or2b_1
X_08673_ _01278_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__nand3_2
XFILLER_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4346__A MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5518_ MuI._1295_ MuI._1297_ MuI._1312_ vssd1 vssd1 vccd1 vccd1 MuI._1313_ sky130_fd_sc_hd__nand3_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07624_ _00131_ _00134_ _00130_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__o21bai_1
XMuI._6498_ MuI._2381_ MuI._2382_ vssd1 vssd1 vccd1 vccd1 MuI._2391_ sky130_fd_sc_hd__nor2_1
XFILLER_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5449_ MuI._1183_ MuI._1235_ MuI._1172_ vssd1 vssd1 vccd1 vccd1 MuI._1237_ sky130_fd_sc_hd__o21a_1
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07555_ _06667_ _06668_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__nand2_1
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10435__A2 _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ _00079_ _00102_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__nor2_1
XFILLER_194_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10386__B _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6212__A2 MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _01810_ _01841_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a21bo_1
XFILLER_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09156_ _01702_ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07976__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__A _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11396__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _00722_ _00723_ _00724_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__and3_1
XFILLER_108_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _01702_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__o21ba_1
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _00653_ _00654_ _00620_ _00655_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__nand4_2
XFILLER_190_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4135__A1_N MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10000_ _01866_ _01867_ _01873_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__nor3_1
XFILLER_89_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _02650_ _02653_ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nor3_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07216__A _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _04547_ _04549_ _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__o211ai_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0915__A1 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _03619_ _03620_ _03634_ _03635_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__nand4_2
XFILLER_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _04683_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__xor2_1
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _03002_ _00002_ _03560_ _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a22o_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4406__D MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4462__A1 MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10764_ _02935_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_201_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _05348_ _05359_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nand2_1
XFILLER_201_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _02707_ _02813_ _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._5411__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695_ _03380_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4422__C MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12179__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12434_ _05269_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__or2_2
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06790__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__B1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__A_N _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _05211_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nand2_1
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5714__A1 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _04082_ _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__and2b_1
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5714__B2 MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _02584_ _04159_ _05021_ _05032_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o311ai_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3725__B1 MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4820_ MuI._0542_ MuI._0543_ vssd1 vssd1 vccd1 vccd1 MuI._0545_ sky130_fd_sc_hd__nor2_1
XFILLER_141_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11247_ _04005_ _04007_ _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a21oi_1
XAuI._1674_ AuI._0119_ AuI._0120_ AuI._0138_ vssd1 vssd1 vccd1 vccd1 AuI._0024_ sky130_fd_sc_hd__or3_1
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._680_ AuI.pe.significand\[2\] AuI.pe.significand\[7\] AuI.pe._197_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._228_ sky130_fd_sc_hd__and3_1
XMuI._4751_ MuI._0466_ MuI._0468_ vssd1 vssd1 vccd1 vccd1 MuI._0469_ sky130_fd_sc_hd__nor2_1
XFILLER_95_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ _03931_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__a21o_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3702_ MuI._2693_ vssd1 vssd1 vccd1 vccd1 MuI._2802_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4682_ MuI._0354_ MuI._0356_ vssd1 vssd1 vccd1 vccd1 MuI._0393_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _02804_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6421_ MuI._2243_ MuI._2305_ vssd1 vssd1 vccd1 vccd1 MuI._2306_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08307__A1 _00596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3633_ MuI.a_operand\[6\] vssd1 vssd1 vccd1 vccd1 MuI._2319_ sky130_fd_sc_hd__clkbuf_4
XFILLER_209_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4166__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6352_ MuI._2228_ MuI._2229_ vssd1 vssd1 vccd1 vccd1 MuI._2230_ sky130_fd_sc_hd__or2b_1
XANTENNA__11871__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3564_ MuI._1538_ MuI._1549_ vssd1 vssd1 vccd1 vccd1 MuI._1560_ sky130_fd_sc_hd__nor2_1
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10665__A2 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__A _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5303_ MuI._3189_ MuI._3190_ MuI.a_operand\[4\] MuI.a_operand\[3\] vssd1 vssd1
+ vccd1 vccd1 MuI._1077_ sky130_fd_sc_hd__and4_1
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6283_ MuI._2145_ MuI._2153_ vssd1 vssd1 vccd1 vccd1 MuI._2155_ sky130_fd_sc_hd__nor2_1
XANTENNA__08883__C _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3495_ MuI._0790_ vssd1 vssd1 vccd1 vccd1 MuI._0801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06684__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5234_ MuI._0932_ MuI._0935_ MuI._0934_ vssd1 vssd1 vccd1 vccd1 MuI._1001_ sky130_fd_sc_hd__o21ba_1
XFILLER_177_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07340_ _06576_ _06577_ _06639_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand4_4
XAuI._1108_ AuI._0262_ AuI._0313_ AuI._0317_ vssd1 vssd1 vccd1 vccd1 AuI._0318_ sky130_fd_sc_hd__a21o_1
XFILLER_177_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5709__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1331__A1 net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5165_ MuI._0921_ MuI._0923_ MuI._0906_ vssd1 vssd1 vccd1 vccd1 MuI._0925_ sky130_fd_sc_hd__a21o_1
X_07271_ _06570_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and2b_1
XAuI._1039_ AuI._0213_ AuI._0250_ vssd1 vssd1 vccd1 vccd1 AuI._0251_ sky130_fd_sc_hd__and2_1
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4116_ MuI._2583_ MuI._2789_ vssd1 vssd1 vccd1 vccd1 MuI._3216_ sky130_fd_sc_hd__nand2_1
XFILLER_164_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09010_ _01537_ _01538_ _01544_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__nand3_1
XANTENNA__07796__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5096_ MuI.a_operand\[12\] MuI.a_operand\[11\] MuI._0017_ MuI._0018_ vssd1 vssd1
+ vccd1 vccd1 MuI._0849_ sky130_fd_sc_hd__and4_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4047_ MuI._3056_ MuI._3126_ MuI._3145_ MuI._3146_ vssd1 vssd1 vccd1 vccd1 MuI._3147_
+ sky130_fd_sc_hd__or4bb_1
XFILLER_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12207__A _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07597__A2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6259__C MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _02522_ _02523_ _02549_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__and3_1
XFILLER_99_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5998_ MuI._1836_ MuI._1840_ MuI._0283_ vssd1 vssd1 vccd1 vccd1 MuI._1841_ sky130_fd_sc_hd__or3b_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12878__B1 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4949_ MuI._0674_ MuI._0678_ MuI._0681_ vssd1 vssd1 vccd1 vccd1 MuI._0687_ sky130_fd_sc_hd__or3_1
XFILLER_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10061__A1_N _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _02248_ _06446_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__nand2_1
XFILLER_101_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _05273_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__and3_1
X_09774_ _02413_ _02421_ _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a21bo_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6619_ MuI._1447_ MuI._1449_ vssd1 vssd1 vccd1 vccd1 MuI._2524_ sky130_fd_sc_hd__nor2_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07036__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08725_ _06515_ _04574_ _00030_ _06519_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__a22o_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4076__A MuI._3158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _01272_ _01273_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__nor2_1
XFILLER_27_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07607_ _00214_ _00223_ _00224_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__nand3_1
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ _01204_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07538_ _06644_ _06645_ _06643_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12802__B1 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1322__A1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07285__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _00081_ _00083_ _00085_ _00086_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08482__B1 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09208_ _01781_ _01780_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10480_ _02959_ _00423_ _05198_ _02905_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a22o_1
XFILLER_136_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10844__B _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _01734_ _01733_ _01732_ _01711_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a211o_1
XANTENNA__12117__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12150_ _04849_ _04941_ _04979_ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a211o_2
XANTENNA__12581__A2 _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11101_ _02759_ _03850_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__nor2_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11956__A _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ _02862_ _05981_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__nand2_1
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12869__B1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09734__B1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11032_ _03774_ _03775_ _03571_ _03741_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__o211a_1
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09426__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11541__B1 _01891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1390_ AuI._0569_ vssd1 vssd1 vccd1 vccd1 AuI._0581_ sky130_fd_sc_hd__inv_2
XFILLER_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6185__B MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3486__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12983_ _05867_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _04702_ _04704_ _04746_ _04748_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a22o_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _04672_ _04673_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__nand3_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816_ _03541_ _03542_ _03537_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a21o_1
X_11796_ _04598_ _04599_ _04426_ _04498_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__o211a_1
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _03416_ _03470_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__xor2_1
XFILLER_158_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12953__C _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ MuI.result\[30\] _02739_ _02745_ _02820_ _06381_ vssd1 vssd1 vccd1 vccd1
+ _06382_ sky130_fd_sc_hd__a221o_1
X_10678_ _03228_ _03282_ _06612_ _04843_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__and4_1
XFILLER_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _05041_ _05151_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__or2_1
XANTENNA__13130__B _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13397_ AuI.result\[28\] _02731_ _06308_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_
+ sky130_fd_sc_hd__a211o_1
XMuI._5921_ MuI._1716_ MuI._1755_ vssd1 vssd1 vccd1 vccd1 MuI._1756_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07766__D net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08776__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12348_ _05191_ _05192_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a21o_1
XFILLER_181_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._801_ AuI.pe._339_ AuI.pe._340_ vssd1 vssd1 vccd1 vccd1 AuI.pe._341_ sky130_fd_sc_hd__nor2b_1
XFILLER_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5852_ MuI._1669_ MuI._1671_ MuI._1678_ vssd1 vssd1 vccd1 vccd1 MuI._1680_ sky130_fd_sc_hd__nand3_1
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10770__A _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ _05037_ _04984_ _05118_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__o211a_2
XANTENNA_AuI.pe._556__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._732_ AuI.pe._062_ AuI.pe._197_ AuI.pe._173_ vssd1 vssd1 vccd1 vccd1 AuI.pe._277_
+ sky130_fd_sc_hd__a21o_1
XMuI._4803_ MuI._0476_ MuI._0490_ MuI._0489_ MuI._0485_ vssd1 vssd1 vccd1 vccd1 MuI._0527_
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5783_ MuI._1598_ MuI._1603_ vssd1 vssd1 vccd1 vccd1 MuI._1605_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1657_ AuI._0008_ AuI._0692_ AuI.operand_a\[27\] AuI._0258_ vssd1 vssd1 vccd1
+ vccd1 AuI._0011_ sky130_fd_sc_hd__a211o_1
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._663_ AuI.pe._211_ AuI.pe._208_ vssd1 vssd1 vccd1 vccd1 AuI.pe._212_ sky130_fd_sc_hd__xor2_1
XMuI._4734_ MuI._0625_ MuI._0246_ MuI._0420_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._0451_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._6112__A1 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _03701_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08597__D _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1588_ AuI._0624_ AuI._0755_ vssd1 vssd1 vccd1 vccd1 AuI._0762_ sky130_fd_sc_hd__or2_1
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._594_ AuI.pe._046_ AuI.pe._112_ AuI.pe._097_ AuI.pe._059_ AuI.pe._147_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._148_ sky130_fd_sc_hd__a221o_1
XMuI._4665_ MuI._0371_ MuI._0373_ MuI._0374_ vssd1 vssd1 vccd1 vccd1 MuI._0375_ sky130_fd_sc_hd__a21bo_1
XFILLER_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06771_ _02959_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__buf_6
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6404_ MuI._2053_ MuI._2085_ MuI._2091_ MuI._2287_ vssd1 vssd1 vccd1 vccd1 MuI._2288_
+ sky130_fd_sc_hd__o31a_1
XMuI._3616_ MuI._1857_ MuI._1879_ MuI._1890_ MuI._2121_ vssd1 vssd1 vccd1 vccd1 MuI._2132_
+ sky130_fd_sc_hd__a31o_1
X_08510_ _00892_ _00893_ _00896_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__nor3_2
XANTENNA_MuI._5862__A2_N MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4596_ MuI._0296_ MuI._0298_ vssd1 vssd1 vccd1 vccd1 MuI._0299_ sky130_fd_sc_hd__nand2_1
X_09490_ _02112_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6335_ MuI._1857_ MuI._1879_ vssd1 vssd1 vccd1 vccd1 MuI._2212_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3547_ MuI._0581_ MuI._0746_ MuI._1164_ MuI._0350_ vssd1 vssd1 vccd1 vccd1 MuI._1373_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08441_ _00858_ _00861_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13037__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6266_ MuI._2134_ MuI._2133_ vssd1 vssd1 vccd1 vccd1 MuI._2136_ sky130_fd_sc_hd__and2b_1
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3478_ MuI._0603_ vssd1 vssd1 vccd1 vccd1 MuI._0614_ sky130_fd_sc_hd__buf_2
X_08372_ _02474_ _06604_ _06580_ _06564_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a22oi_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5217_ MuI._0952_ MuI._0953_ MuI._0975_ MuI._0981_ vssd1 vssd1 vccd1 vccd1 MuI._0982_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07323_ _06585_ _06622_ _06623_ _06517_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and4_1
XFILLER_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6197_ MuI._2594_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._2060_ sky130_fd_sc_hd__nand2_1
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5148_ MuI._0871_ MuI._0880_ MuI._0879_ vssd1 vssd1 vccd1 vccd1 MuI._0906_ sky130_fd_sc_hd__a21bo_1
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07254_ _06542_ _06543_ _06552_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a21o_1
XFILLER_165_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5079_ MuI._2845_ MuI._0110_ MuI._0244_ MuI._2844_ vssd1 vssd1 vccd1 vccd1 MuI._0830_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07185_ _06470_ _06467_ _06468_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__or3_1
XANTENNA__08134__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08767__A1 _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12563__A2 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B2 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10680__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12315__A2 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__B _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3703__A MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09826_ _02469_ _02477_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand3_2
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ _02387_ _02389_ _02380_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06969_ net14 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__buf_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _01323_ _01325_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__xnor2_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09688_ _02328_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__nor2_1
XANTENNA__11826__B2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4417__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _01249_ _01251_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13028__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4417__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11016__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07213__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ _04440_ _04442_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__xor2_4
XANTENNA_MuI._5349__B MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _02752_ _03129_ _03130_ _03313_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__a31o_2
XANTENNA__07258__A1 _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _02658_ net39 _03082_ _00789_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__and4_1
XANTENNA__08455__B1 _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10262__B1 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ _03236_ _03237_ _03221_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__a21o_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _06227_ _06172_ _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__o21a_1
XFILLER_155_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _02834_ _06096_ _02836_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a21oi_1
X_10463_ _03159_ _03162_ _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__nand3_2
XFILLER_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._0890_ net57 net129 vssd1 vssd1 vccd1 vccd1 AuI._0110_ sky130_fd_sc_hd__xnor2_4
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08758__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _04810_ _04938_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nor2_1
XANTENNA__08758__B2 _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ _02687_ _02688_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__nor2_1
XFILLER_182_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input67_A b_operand[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__or2_1
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12133_ _00292_ _00002_ _04960_ _04962_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__a22o_1
XANTENNA_AuI._0828__B net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1511_ AuI.operand_a\[28\] AuI.operand_a\[29\] AuI._0604_ vssd1 vssd1 vccd1 vccd1
+ AuI._0697_ sky130_fd_sc_hd__nand3_1
X_12064_ MuI.result\[12\] _02739_ _04886_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09156__A _01702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08060__A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4709__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12711__C1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _03757_ _03758_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__nor2_1
XFILLER_49_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1442_ AuI._0623_ AuI._0624_ AuI._0625_ AuI._0626_ AuI._0627_ vssd1 vssd1 vccd1
+ vccd1 AuI._0628_ sky130_fd_sc_hd__o2111a_1
XANTENNA__10868__A2 _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07733__A2 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1373_ AuI._0559_ AuI._0564_ vssd1 vssd1 vccd1 vccd1 AuI._0565_ sky130_fd_sc_hd__xor2_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4450_ MuI._0131_ MuI._0136_ MuI._0137_ vssd1 vssd1 vccd1 vccd1 MuI._0138_ sky130_fd_sc_hd__a21o_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _02751_ _05774_ _05775_ _05857_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__a31o_4
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4381_ MuI._0060_ MuI._0062_ vssd1 vssd1 vccd1 vccd1 MuI._0063_ sky130_fd_sc_hd__nand2_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _04728_ _04729_ _04724_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__a21o_1
XANTENNA__13125__B _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11293__A2 _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6120_ MuI._1971_ MuI._1974_ vssd1 vssd1 vccd1 vccd1 MuI._1975_ sky130_fd_sc_hd__xnor2_4
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12897_ _03346_ _05906_ _05981_ _03293_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a22o_1
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _00878_ _03444_ _05948_ _00012_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a22o_1
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4163__B MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6051_ MuI._1893_ MuI._1898_ vssd1 vssd1 vccd1 vccd1 MuI._1899_ sky130_fd_sc_hd__xor2_1
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6081__D MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07249__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5002_ MuI._0552_ MuI._0554_ MuI._0553_ vssd1 vssd1 vccd1 vccd1 MuI._0745_ sky130_fd_sc_hd__o21ai_1
X_11779_ _04579_ _04580_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
XFILLER_202_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10253__B1 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08235__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13449_ _02820_ _02821_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__or2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08749__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08749__B2 _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5904_ MuI._0750_ MuI._1685_ MuI._1686_ MuI._1696_ vssd1 vssd1 vccd1 vccd1 MuI._1738_
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07421__A1 _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__B _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07421__B2 _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08990_ _01605_ _01606_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__nand3_1
XFILLER_69_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5835_ MuI._1558_ MuI._1564_ MuI._1661_ vssd1 vssd1 vccd1 vccd1 MuI._1662_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09066__A _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _00554_ _00558_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__and2_1
XAuI.pe._715_ AuI.pe._145_ AuI.pe._096_ AuI.pe._118_ AuI.pe._380_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._261_ sky130_fd_sc_hd__a22o_1
XANTENNA__12204__B _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08401__C _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5766_ MuI._2803_ MuI._2829_ MuI._3246_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._1586_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_205_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07872_ _00283_ _04251_ _00487_ _00488_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__nand4_2
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6097__B1 MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._646_ AuI.pe._063_ AuI.pe._133_ AuI.pe._173_ AuI.pe._055_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._196_ sky130_fd_sc_hd__a22o_1
XMuI._4717_ MuI._0430_ MuI._0431_ MuI._2473_ MuI._3372_ vssd1 vssd1 vccd1 vccd1 MuI._0432_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09611_ _02118_ _02205_ _04358_ _00083_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__nand4_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5697_ MuI._1507_ MuI._1508_ MuI._1509_ vssd1 vssd1 vccd1 vccd1 MuI._1510_ sky130_fd_sc_hd__nand3b_1
X_06823_ _03518_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._577_ AuI.pe.significand\[12\] AuI.pe._388_ AuI.pe._389_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._132_ sky130_fd_sc_hd__and3_1
XMuI._4648_ MuI._0349_ MuI._0355_ vssd1 vssd1 vccd1 vccd1 MuI._0356_ sky130_fd_sc_hd__and2_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06754_ _02776_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[12\] sky130_fd_sc_hd__clkbuf_1
X_09542_ _06545_ _04251_ _02171_ _02172_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a31o_1
XANTENNA__12220__A _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4579_ MuI._0277_ MuI._0279_ vssd1 vssd1 vccd1 vccd1 MuI._0280_ sky130_fd_sc_hd__or2b_1
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06685_ _02031_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__buf_2
X_09473_ _06491_ _04509_ _00035_ _06534_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a22oi_2
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3870__A2 MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6318_ MuI._2191_ MuI._2192_ vssd1 vssd1 vccd1 vccd1 MuI._2193_ sky130_fd_sc_hd__nor2_1
XFILLER_197_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _01040_ _01041_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__nor2_1
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5072__A1 MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._441__A AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6249_ MuI._2115_ MuI._2116_ vssd1 vssd1 vccd1 vccd1 MuI._2117_ sky130_fd_sc_hd__and2_1
X_08355_ _06488_ _06517_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__nand2_1
XFILLER_165_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07306_ _06601_ _06603_ _06605_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08790__D _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ _00873_ _00872_ _00871_ _00849_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__a211o_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07237_ _02205_ _06537_ _05756_ _02118_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__a22oi_4
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12536__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11002__C _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ net37 vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__buf_4
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07099_ _05209_ _06284_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__and2_1
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__B1 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09126__D _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _00150_ net126 net125 _06469_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XFILLER_19_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11953__B _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12820_ _00292_ _05649_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__nand2_2
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07224__A _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12751_ _05535_ _05539_ _05624_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a211o_1
XFILLER_54_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _04383_ _04422_ _04423_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__nor3_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05511_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nor3_2
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6260__B1 MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _04422_ _04423_ _04383_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__o21ai_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11564_ _02790_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__xor2_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__A2 _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _05671_ _02727_ _04627_ FuI.Integer\[26\] vssd1 vssd1 vccd1 vccd1 _06214_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10515_ _03069_ _03077_ _03076_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a21o_1
XAuI._0942_ AuI._0113_ AuI._0118_ vssd1 vssd1 vccd1 vccd1 AuI._0154_ sky130_fd_sc_hd__nand2_2
XANTENNA__07651__A1 _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _02987_ _04854_ _04274_ _04275_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__nand4_1
XANTENNA__07651__B2 _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4963__A2_N MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10446_ _02965_ _04251_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__nand2_1
X_13234_ _06139_ _06141_ _06142_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0873_ AuI._0086_ AuI._0090_ AuI._0092_ vssd1 vssd1 vccd1 vccd1 AuI._0093_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10538__A1 _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10538__B2 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3950_ MuI._2055_ MuI._2693_ MuI._2918_ MuI._1472_ vssd1 vssd1 vccd1 vccd1 MuI._3050_
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _02431_ _02485_ _00382_ _00163_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__nand4_1
X_13165_ _06066_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__nand2_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__C _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3881_ MuI._2978_ MuI._2979_ MuI._2980_ vssd1 vssd1 vccd1 vccd1 MuI._2981_ sky130_fd_sc_hd__nand3_1
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _00534_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a21bo_1
X_13096_ _02782_ _05995_ _02713_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5620_ MuI._1382_ MuI._1424_ vssd1 vssd1 vccd1 vccd1 MuI._1425_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _04755_ _04757_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__nor2_1
XAuI.pe._500_ AuI.pe._020_ AuI.pe._054_ AuI.pe._058_ AuI.pe._061_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[4\] sky130_fd_sc_hd__a211o_1
XANTENNA__07167__B1 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5551_ MuI._1308_ MuI._1306_ MuI._1305_ vssd1 vssd1 vccd1 vccd1 MuI._1349_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1425_ AuI._0609_ AuI._0610_ vssd1 vssd1 vccd1 vccd1 AuI._0611_ sky130_fd_sc_hd__and2b_1
XAuI.pe._431_ AuI.pe._392_ AuI.pe._397_ vssd1 vssd1 vccd1 vccd1 AuI.pe._398_ sky130_fd_sc_hd__nor2_1
XMuI._4502_ MuI._0192_ MuI._0194_ vssd1 vssd1 vccd1 vccd1 MuI._0195_ sky130_fd_sc_hd__nand2_1
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5482_ MuI._1261_ MuI._1264_ vssd1 vssd1 vccd1 vccd1 MuI._1273_ sky130_fd_sc_hd__and2_1
XAuI._1356_ net14 net46 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0550_ sky130_fd_sc_hd__mux2_2
XFILLER_92_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4433_ MuI._0094_ MuI._0118_ vssd1 vssd1 vccd1 vccd1 MuI._0120_ sky130_fd_sc_hd__nor2_1
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09052__C _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1287_ AuI._0420_ AuI._0465_ AuI._0474_ vssd1 vssd1 vccd1 vccd1 AuI._0486_ sky130_fd_sc_hd__and3_1
XANTENNA__11266__A2 _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _05748_ _05752_ _05746_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21boi_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4364_ MuI._3316_ MuI._0044_ vssd1 vssd1 vccd1 vccd1 MuI._0045_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5054__A1 MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6103_ MuI._1941_ MuI._1955_ vssd1 vssd1 vccd1 vccd1 MuI._1957_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._5054__B2 MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4295_ MuI._3312_ MuI._3394_ vssd1 vssd1 vccd1 vccd1 MuI._3395_ sky130_fd_sc_hd__nor2_1
XANTENNA__11018__A2 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4902__A MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6034_ MuI._1850_ MuI._1880_ vssd1 vssd1 vccd1 vccd1 MuI._1881_ sky130_fd_sc_hd__xor2_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08140_ net122 _06562_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__nand2_1
XFILLER_193_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08071_ _00687_ _00688_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__nor2_2
XFILLER_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _05660_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6306__A1 MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__A2_N _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08412__B _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6857__A2 MuI._2733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07309__A _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6867_ MuI._2768_ MuI._2493_ vssd1 vssd1 vccd1 vccd1 MuI._2769_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08973_ _01566_ _01567_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA_MuI._4349__A MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5818_ MuI._1462_ MuI._1555_ vssd1 vssd1 vccd1 vccd1 MuI._1643_ sky130_fd_sc_hd__nand2_1
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6798_ MuI._2685_ MuI._2596_ MuI._2600_ MuI._2612_ vssd1 vssd1 vccd1 vccd1 MuI._2721_
+ sky130_fd_sc_hd__or4_1
X_07924_ _00533_ _00541_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5749_ MuI._1467_ MuI._1469_ MuI._1566_ vssd1 vssd1 vccd1 vccd1 MuI._1567_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11773__B _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _00455_ _00456_ _00471_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__o21a_1
XFILLER_84_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._629_ AuI.pe._145_ AuI.pe._041_ AuI.pe._078_ AuI.pe._393_ AuI.pe._180_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._181_ sky130_fd_sc_hd__a221o_1
XANTENNA__13046__A _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ _03335_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__buf_4
X_07786_ _00402_ _00403_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__and2b_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07044__A _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _01999_ _02061_ _02067_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__or3_1
XFILLER_37_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06737_ _02593_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__buf_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _02077_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__nor2_1
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06883__A _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _02582_ _02647_ _00032_ _04767_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__and4_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._111_ FuI.a_operand\[26\] FuI._037_ vssd1 vssd1 vccd1 vccd1 FuI._023_ sky130_fd_sc_hd__or2b_1
X_09387_ _02851_ _03884_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nand2_1
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ _00817_ _00954_ _00818_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__and3_1
XANTENNA__10110__A_N _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10768__B2 _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _00883_ _00886_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._5346__C MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4250__C MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ _02986_ _02988_ _02979_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a21o_1
XFILLER_165_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12509__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _04041_ _04042_ _04033_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__a21o_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ _02876_ _02910_ _02914_ _02829_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a211oi_4
XFILLER_180_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11193__A1 _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5362__B MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _02838_ _02839_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nor2_2
XANTENNA__07219__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10940__A1 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10940__B2 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5520__A2 MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _02259_ _04057_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12693__A1 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08897__B1 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._1210_ net34 net66 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0415_ sky130_fd_sc_hd__mux2_2
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08361__A2 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09153__B _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4087__A2 MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1141_ AuI._0329_ AuI._0349_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[3\]
+ sky130_fd_sc_hd__xnor2_4
X_12803_ _05598_ _05670_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or3_4
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _03734_ _03735_ _03591_ _03594_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__a211o_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _03174_ _05970_ _05496_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__and3_1
XAuI._1072_ AuI._0199_ AuI._0200_ AuI._0282_ AuI._0205_ vssd1 vssd1 vccd1 vccd1 AuI._0283_
+ sky130_fd_sc_hd__a31o_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12665_ _05529_ _05533_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand3_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3598__A1 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3598__B2 MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4080_ MuI._3157_ MuI._3179_ vssd1 vssd1 vccd1 vccd1 MuI._3180_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11204__A _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11616_ _00086_ _00081_ _06476_ _06489_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and4_1
XFILLER_168_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12596_ _05458_ _05459_ _05440_ _05322_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__o211ai_1
XFILLER_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _02550_ _02724_ _04329_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a211o_1
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output98_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0925_ AuI._0116_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[30\] sky130_fd_sc_hd__inv_2
XANTENNA__11858__B _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11478_ _02965_ _04660_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nand2_1
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4982_ MuI._0626_ MuI._0628_ vssd1 vssd1 vccd1 vccd1 MuI._0723_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13173__A2 _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ _06107_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__xor2_1
X_10429_ _02767_ _02882_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__xnor2_1
XAuI._0856_ AuI._0070_ net40 net122 AuI._0074_ AuI._0075_ vssd1 vssd1 vccd1 vccd1
+ AuI._0076_ sky130_fd_sc_hd__a221oi_1
XFILLER_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3933_ MuI._3027_ MuI._3031_ MuI._3032_ vssd1 vssd1 vccd1 vccd1 MuI._3033_ sky130_fd_sc_hd__o21ba_1
XFILLER_140_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6721_ MuI._2629_ MuI._2635_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2636_ sky130_fd_sc_hd__mux2_1
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10481__C _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05980_ _05979_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__and2b_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4169__A MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6652_ MuI._1829_ MuI._2512_ vssd1 vssd1 vccd1 vccd1 MuI._2560_ sky130_fd_sc_hd__or2b_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3864_ MuI._2961_ MuI._2962_ MuI._2963_ vssd1 vssd1 vccd1 vccd1 MuI._2964_ sky130_fd_sc_hd__nand3b_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11874__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _05881_ _05899_ _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__o21ai_1
XMuI._5603_ MuI._1292_ MuI._1293_ MuI._1404_ vssd1 vssd1 vccd1 vccd1 MuI._1407_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6583_ MuI._0999_ MuI._2482_ MuI._2483_ vssd1 vssd1 vccd1 vccd1 MuI._2485_ sky130_fd_sc_hd__or3_2
XMuI._3795_ MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 MuI._2895_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5534_ MuI._1287_ MuI._1291_ MuI._1294_ MuI._1330_ vssd1 vssd1 vccd1 vccd1 MuI._1331_
+ sky130_fd_sc_hd__nand4_2
XAuI._1408_ AuI._0576_ AuI._0583_ vssd1 vssd1 vccd1 vccd1 AuI._0597_ sky130_fd_sc_hd__nor2_1
XANTENNA__09063__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07640_ _03099_ _04358_ _04445_ _03056_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__a22oi_1
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._414_ AuI.pe._378_ AuI.pe._379_ AuI.pe._380_ vssd1 vssd1 vccd1 vccd1 AuI.pe._381_
+ sky130_fd_sc_hd__or3b_1
XFILLER_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5465_ MuI.a_operand\[6\] MuI.a_operand\[5\] MuI._3262_ MuI._0020_ vssd1 vssd1
+ vccd1 vccd1 MuI._1255_ sky130_fd_sc_hd__and4_1
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1339_ AuI._0528_ AuI._0534_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[16\]
+ sky130_fd_sc_hd__xor2_1
X_07571_ _06680_ _06525_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__nand2_1
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4416_ MuI._0100_ vssd1 vssd1 vccd1 vccd1 MuI._0101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09310_ _01927_ _01886_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__xnor2_1
XMuI._5396_ MuI._1176_ MuI._1177_ vssd1 vssd1 vccd1 vccd1 MuI._1179_ sky130_fd_sc_hd__nand2_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4347_ MuI._0025_ MuI._3399_ vssd1 vssd1 vccd1 vccd1 MuI._0026_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _01262_ _01264_ _01266_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__nor3_1
XFILLER_210_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3589__A1 MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08407__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4278_ MuI._3357_ MuI._3358_ MuI._3377_ vssd1 vssd1 vccd1 vccd1 MuI._3378_ sky130_fd_sc_hd__nor3_1
X_09172_ _01717_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a21o_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4351__B MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6017_ MuI._1860_ MuI._1861_ vssd1 vssd1 vccd1 vccd1 MuI._1862_ sky130_fd_sc_hd__xor2_1
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _00737_ _00738_ _00739_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__a21o_1
XANTENNA__11947__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07615__A1 _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08054_ _00670_ _00518_ _00671_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a21boi_4
XFILLER_190_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07005_ _05478_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[23\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_MuI._5463__A MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07039__A _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5613__D MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08956_ _01571_ _01573_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06878__A _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0926__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4710__B1 MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07907_ _00366_ _00368_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__or2b_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _01497_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__xor2_1
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09540__A1 _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09540__B2 _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07838_ _00452_ _00453_ _00454_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__a21oi_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07769_ _00384_ _00386_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__nor2_1
XFILLER_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09508_ _02127_ _02128_ _02135_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__and3_1
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10780_ _02769_ _02770_ _02928_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a21o_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09439_ _06680_ _04035_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__o2bb2a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _05301_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__nand2_1
XFILLER_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4261__B MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _02887_ _02759_ _03850_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o31ai_1
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12381_ _05114_ _05145_ _05228_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__o211ai_4
XFILLER_138_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ _04725_ _04098_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ _03945_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__inv_2
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11166__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__B2 _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13002_ _05882_ _05811_ _05893_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and3_1
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ _02845_ _02896_ _02846_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a21oi_1
X_11194_ _00444_ _05327_ _03949_ _03950_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__nand4_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10145_ _05853_ _03680_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and2b_1
XFILLER_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06788__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12115__B1 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4139__D MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _06428_ _02704_ _02716_ _02748_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__o211ai_4
XFILLER_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6635__C MuI._2534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3580_ MuI._0988_ MuI._1725_ vssd1 vssd1 vccd1 vccd1 MuI._1736_ sky130_fd_sc_hd__nand2_1
XANTENNA__10677__B1 _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5257__A1 MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5250_ MuI.b_operand\[8\] MuI._0088_ vssd1 vssd1 vccd1 vccd1 MuI._1018_ sky130_fd_sc_hd__nand2_1
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1124_ AuI._0330_ AuI._0331_ AuI._0332_ vssd1 vssd1 vccd1 vccd1 AuI._0333_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09611__B _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4201_ MuI._3298_ MuI._3300_ vssd1 vssd1 vccd1 vccd1 MuI._3301_ sky130_fd_sc_hd__or2b_1
XFILLER_16_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _00281_ _03443_ _00040_ _04789_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nand4_1
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5181_ MuI._2803_ MuI._0110_ MuI._0244_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._0942_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07412__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12717_ _03489_ _05582_ _05583_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a31o_1
XANTENNA__07845__A1 _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1055_ AuI._0199_ AuI._0200_ AuI._0224_ vssd1 vssd1 vccd1 vccd1 AuI._0266_ sky130_fd_sc_hd__and3_1
XANTENNA__07845__B2 _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4132_ MuI._3230_ MuI._3231_ vssd1 vssd1 vccd1 vccd1 MuI._3232_ sky130_fd_sc_hd__or2_1
XFILLER_176_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12648_ _06439_ _05327_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__nand2_1
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4063_ MuI._2887_ MuI._3162_ MuI._2968_ vssd1 vssd1 vccd1 vccd1 MuI._3163_ sky130_fd_sc_hd__a21o_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _05310_ _05318_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0908_ AuI._0127_ vssd1 vssd1 vccd1 vccd1 AuI.exp_a sky130_fd_sc_hd__buf_2
XFILLER_171_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._141__147 vssd1 vssd1 vccd1 vccd1 FuI._141__147/HI net147 sky130_fd_sc_hd__conb_1
XANTENNA_MuI._6098__B MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4965_ MuI._0701_ MuI._0704_ vssd1 vssd1 vccd1 vccd1 MuI._0705_ sky130_fd_sc_hd__and2_1
XFILLER_171_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0839_ net115 net37 vssd1 vssd1 vccd1 vccd1 AuI._0059_ sky130_fd_sc_hd__and2b_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6704_ MuI._2384_ MuI._2603_ MuI._2392_ vssd1 vssd1 vccd1 vccd1 MuI._2618_ sky130_fd_sc_hd__o21ai_2
XMuI._3916_ MuI._0867_ MuI._2791_ vssd1 vssd1 vccd1 vccd1 MuI._3016_ sky130_fd_sc_hd__nand2_1
X_08810_ _01419_ _01422_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__xnor2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4896_ MuI._0626_ MuI._0628_ vssd1 vssd1 vccd1 vccd1 MuI._0629_ sky130_fd_sc_hd__nand2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _02376_ _02383_ _02382_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o21ai_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6635_ MuI._2514_ MuI._2518_ MuI._2534_ MuI._2541_ vssd1 vssd1 vccd1 vccd1 MuI._2542_
+ sky130_fd_sc_hd__or4_1
XMuI._3847_ MuI._2330_ MuI._0438_ vssd1 vssd1 vccd1 vccd1 MuI._2947_ sky130_fd_sc_hd__nand2_1
XFILLER_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _06598_ _06599_ _04294_ _00072_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__and4_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6566_ MuI._2464_ MuI._2465_ vssd1 vssd1 vccd1 vccd1 MuI._2466_ sky130_fd_sc_hd__or2_1
XFILLER_66_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3778_ MuI._2870_ MuI._2872_ MuI._2877_ vssd1 vssd1 vccd1 vccd1 MuI._2878_ sky130_fd_sc_hd__or3_1
X_08672_ _00983_ _00977_ _00982_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4346__B MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5517_ MuI._1302_ MuI._1310_ MuI._1311_ vssd1 vssd1 vccd1 vccd1 MuI._1312_ sky130_fd_sc_hd__a21bo_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6497_ MuI._2240_ MuI._2389_ MuI._2239_ vssd1 vssd1 vccd1 vccd1 MuI._2390_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12409__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _00238_ _00239_ _00236_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__a21o_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5448_ MuI._1178_ MuI._1183_ MuI._1235_ vssd1 vssd1 vccd1 vccd1 MuI._1236_ sky130_fd_sc_hd__nor3_2
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07554_ _00168_ _00170_ _00169_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__a21o_1
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07322__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5379_ MuI._1063_ MuI._1066_ vssd1 vssd1 vccd1 vccd1 MuI._1160_ sky130_fd_sc_hd__xnor2_1
XFILLER_210_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07485_ _00079_ _00102_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__and2_1
XFILLER_195_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10386__C _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ _01837_ _01840_ _01811_ _01758_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o211ai_1
XFILLER_107_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _01704_ _01703_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nor2_1
XANTENNA__07976__B _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10683__A _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A1 _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__B2 AuI.result\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08106_ _00442_ _00451_ _00450_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a21bo_1
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ _02420_ _06513_ _00084_ _04574_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__and4_1
XFILLER_163_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _00588_ _00619_ _00614_ _00618_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__o211ai_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _02649_ _02648_ _01865_ _02646_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o211a_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__A1_N _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08939_ _02851_ _04380_ _01246_ _01247_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11019__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _02752_ _04637_ _04639_ _04765_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__a31o_4
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07524__B1 _00141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._624__A AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _03619_ _03620_ _03634_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a22o_1
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ _04690_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__and2b_1
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10832_ _00049_ _00046_ _05252_ _00412_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nand4_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13073__A1 _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4462__A2 MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11084__B1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5368__A MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4272__A MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10763_ _03329_ _03485_ _03133_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o21a_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _05348_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__or2_1
XANTENNA__10831__B1 _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5411__A1 MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ _02705_ _02812_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__nand2_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10694_ _03412_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__nand2_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5411__B2 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4422__D MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _05275_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09159__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12364_ _03733_ _05047_ _05210_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21o_1
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08063__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _04078_ _04080_ _04081_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__a21o_1
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5714__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ _05136_ _06427_ _05137_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or3b_1
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1673_ AuI._0116_ AuI._0695_ AuI._0021_ AuI._0023_ vssd1 vssd1 vccd1 vccd1 AuI.result\[30\]
+ sky130_fd_sc_hd__a31oi_1
X_11246_ _03133_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__nand2_1
XFILLER_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12887__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0847__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4750_ MuI._0466_ MuI._0467_ MuI._2451_ MuI.b_operand\[8\] vssd1 vssd1 vccd1
+ vccd1 MuI._0468_ sky130_fd_sc_hd__and4bb_1
XFILLER_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13409__A _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10197__B_N _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _03931_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand3_1
XMuI._3701_ MuI._2649_ MuI._2682_ MuI._2528_ MuI._2800_ vssd1 vssd1 vccd1 vccd1 MuI._2801_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07939__A1_N _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4681_ MuI._0385_ MuI._0389_ MuI._0391_ vssd1 vssd1 vccd1 vccd1 MuI._0392_ sky130_fd_sc_hd__or3_1
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _02802_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nor2_1
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6420_ MuI._2300_ MuI._2304_ vssd1 vssd1 vccd1 vccd1 MuI._2305_ sky130_fd_sc_hd__nor2_1
XMuI._3632_ MuI._1758_ MuI._2297_ vssd1 vssd1 vccd1 vccd1 MuI._2308_ sky130_fd_sc_hd__nor2_1
XANTENNA__09504__A1 _01891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A2 _00919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10059_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__buf_2
XFILLER_208_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._740__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4166__B MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6351_ MuI._2208_ MuI._2210_ MuI._2227_ vssd1 vssd1 vccd1 vccd1 MuI._2229_ sky130_fd_sc_hd__or3b_1
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3563_ MuI._1109_ MuI._1252_ vssd1 vssd1 vccd1 vccd1 MuI._1549_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11871__B _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5302_ MuI._3190_ MuI.a_operand\[4\] MuI._0304_ MuI._3189_ vssd1 vssd1 vccd1
+ vccd1 MuI._1075_ sky130_fd_sc_hd__a22o_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6282_ MuI._2151_ MuI._2152_ vssd1 vssd1 vccd1 vccd1 MuI._2153_ sky130_fd_sc_hd__nor2_1
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3494_ MuI._0779_ vssd1 vssd1 vccd1 vccd1 MuI._0790_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08883__D _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5233_ MuI._0995_ MuI._0998_ vssd1 vssd1 vccd1 vccd1 MuI._1000_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1107_ AuI._0152_ AuI._0236_ AuI._0316_ AuI._0246_ vssd1 vssd1 vccd1 vccd1 AuI._0317_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07142__A _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5164_ MuI._0906_ MuI._0921_ MuI._0923_ vssd1 vssd1 vccd1 vccd1 MuI._0924_ sky130_fd_sc_hd__nand3_2
XFILLER_177_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ _06567_ _06569_ _06559_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a21o_1
XAuI._1038_ AuI._0235_ AuI._0247_ AuI._0249_ vssd1 vssd1 vccd1 vccd1 AuI._0250_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4115_ MuI._3212_ MuI._3214_ vssd1 vssd1 vccd1 vccd1 MuI._3215_ sky130_fd_sc_hd__xnor2_1
XMuI._5095_ MuI._2765_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0848_ sky130_fd_sc_hd__nand2_1
XANTENNA__11599__A _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4046_ MuI._3142_ MuI._3143_ MuI._3144_ vssd1 vssd1 vccd1 vccd1 MuI._3146_ sky130_fd_sc_hd__a21o_1
XFILLER_145_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12207__B _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._559__B1 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09911_ _02548_ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__and2_1
XANTENNA_AuI.pe._709__A AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5997_ MuI._0551_ MuI._1837_ MuI._1839_ vssd1 vssd1 vccd1 vccd1 MuI._1840_ sky130_fd_sc_hd__nand3_1
XANTENNA__12878__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4948_ MuI._0683_ MuI._0685_ vssd1 vssd1 vccd1 vccd1 MuI._0686_ sky130_fd_sc_hd__nor2_1
X_09842_ _02493_ _02495_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11550__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4879_ MuI._0607_ MuI._0608_ MuI._0598_ MuI._0602_ vssd1 vssd1 vccd1 vccd1 MuI._0610_
+ sky130_fd_sc_hd__a211o_1
X_09773_ _02414_ _02415_ _02419_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nand3_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3899__C MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06985_ _05262_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__clkbuf_4
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6618_ MuI._1447_ MuI._1449_ vssd1 vssd1 vccd1 vccd1 MuI._2523_ sky130_fd_sc_hd__and2_1
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08724_ _01336_ _01341_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__or2b_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6549_ MuI._2434_ MuI._2436_ vssd1 vssd1 vccd1 vccd1 MuI._2447_ sky130_fd_sc_hd__nor2_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08655_ _01245_ _01269_ _01271_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__nor3_1
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10678__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _00220_ _00222_ _00215_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a21o_1
XFILLER_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08586_ _00095_ _00096_ _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__and4_1
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07052__A _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07537_ _00151_ _00152_ _00154_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__or3_1
XANTENNA__12802__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4523__C MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07987__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06891__A _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07285__A2 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ net118 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__buf_4
XANTENNA__08482__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08482__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ _01812_ _01823_ _01824_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__nand3_2
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ _00007_ _00008_ _00015_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21o_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10844__C _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _01753_ _01754_ _01747_ _01750_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__o211a_1
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5635__B MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__B _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5157__B1 MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ _01596_ _01595_ _01594_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__o21ai_1
XFILLER_151_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _03683_ _03685_ _02758_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09707__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ _04856_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__inv_2
XANTENNA__11956__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08611__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11031_ _03571_ _03741_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a211oi_4
XANTENNA__09426__B _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6185__C MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _05872_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A a_operand[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _04702_ _04704_ _04746_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__nand4_2
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _04518_ _04523_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nand2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _03537_ _03541_ _03542_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nand3_2
XFILLER_60_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _04426_ _04498_ _04598_ _04599_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a211oi_1
XFILLER_201_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10746_ _03467_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5826__A MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ _05917_ _02728_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__nor2_1
XFILLER_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10677_ _00727_ _04789_ _00445_ _00728_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12308__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ _05149_ _05157_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ MuI.result\[28\] _02736_ _02944_ _05724_ _06309_ vssd1 vssd1 vccd1 vccd1
+ _06310_ sky130_fd_sc_hd__a221o_1
XFILLER_154_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5920_ MuI._1717_ MuI._1754_ vssd1 vssd1 vccd1 vccd1 MuI._1755_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08224__C _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A2 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _05096_ _05098_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__nand2_1
XFILLER_181_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._800_ AuI.pe._331_ AuI.pe._333_ AuI.pe._338_ AuI.operand_a\[25\] vssd1 vssd1
+ vccd1 vccd1 AuI.pe._340_ sky130_fd_sc_hd__a31o_1
XFILLER_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12309__B1 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output80_A net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5851_ MuI._1669_ MuI._1671_ MuI._1678_ vssd1 vssd1 vccd1 vccd1 MuI._1679_ sky130_fd_sc_hd__a21o_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _05116_ _05117_ _05075_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a21o_1
XANTENNA__08521__A _01096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._731_ AuI.pe._020_ AuI.pe._274_ AuI.pe._275_ vssd1 vssd1 vccd1 vccd1 AuI.pe._276_
+ sky130_fd_sc_hd__a21o_1
XMuI._4802_ MuI._0521_ MuI._0522_ MuI._0517_ MuI._0520_ vssd1 vssd1 vccd1 vccd1 MuI._0525_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5782_ MuI._1599_ MuI._1602_ vssd1 vssd1 vccd1 vccd1 MuI._1603_ sky130_fd_sc_hd__xnor2_1
X_11229_ _03987_ _03988_ _03812_ _03815_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__o211ai_2
XFILLER_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1656_ AuI._0010_ vssd1 vssd1 vccd1 vccd1 AuI.result\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._662_ AuI.pe.significand\[17\] vssd1 vssd1 vccd1 vccd1 AuI.pe._211_ sky130_fd_sc_hd__buf_2
XMuI._4733_ MuI._0443_ MuI._0448_ vssd1 vssd1 vccd1 vccd1 MuI._0450_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6112__A2 MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1587_ AuI._0630_ AuI._0623_ vssd1 vssd1 vccd1 vccd1 AuI._0761_ sky130_fd_sc_hd__or2_1
XANTENNA__12978__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4664_ MuI._0236_ MuI._0249_ MuI._0369_ vssd1 vssd1 vccd1 vccd1 MuI._0374_ sky130_fd_sc_hd__o21ai_1
XAuI.pe._593_ AuI.pe._072_ AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 AuI.pe._147_ sky130_fd_sc_hd__and2_1
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06770_ _02948_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__buf_6
XANTENNA__06976__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6403_ MuI._2092_ MuI._2097_ vssd1 vssd1 vccd1 vccd1 MuI._2287_ sky130_fd_sc_hd__nand2_1
XMuI._3615_ MuI._1912_ MuI._2110_ vssd1 vssd1 vccd1 vccd1 MuI._2121_ sky130_fd_sc_hd__nor2_1
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4595_ MuI._0289_ MuI._0297_ vssd1 vssd1 vccd1 vccd1 MuI._0298_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6334_ MuI._2163_ MuI._2166_ vssd1 vssd1 vccd1 vccd1 MuI._2211_ sky130_fd_sc_hd__or2b_1
XMuI._3546_ MuI._1208_ MuI._1351_ vssd1 vssd1 vccd1 vccd1 MuI._1362_ sky130_fd_sc_hd__or2_1
XFILLER_63_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _01009_ _01013_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__or2b_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13037__B2 _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6265_ MuI._2133_ MuI._2134_ vssd1 vssd1 vccd1 vccd1 MuI._2135_ sky130_fd_sc_hd__and2b_1
XMuI._3477_ MuI.b_operand\[21\] vssd1 vssd1 vccd1 vccd1 MuI._0603_ sky130_fd_sc_hd__buf_2
X_08371_ net106 _06602_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__nand2_1
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10212__B_N _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5216_ MuI._0978_ MuI._0980_ vssd1 vssd1 vccd1 vccd1 MuI._0981_ sky130_fd_sc_hd__or2_1
XMuI._6196_ MuI._2057_ MuI._2058_ vssd1 vssd1 vccd1 vccd1 MuI._2059_ sky130_fd_sc_hd__nor2_1
X_07322_ net14 vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__clkbuf_8
XFILLER_177_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08464__A1 _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5147_ MuI._0903_ MuI._0904_ vssd1 vssd1 vccd1 vccd1 MuI._0905_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1347__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ _06474_ _06484_ _06473_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__a21bo_1
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12218__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5078_ MuI._2836_ MuI._2838_ MuI._0444_ MuI.a_operand\[1\] vssd1 vssd1 vccd1
+ vccd1 MuI._0829_ sky130_fd_sc_hd__and4_1
XFuI._147__153 vssd1 vssd1 vccd1 vccd1 FuI._147__153/HI net153 sky130_fd_sc_hd__conb_1
X_07184_ _06473_ _06474_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nand3_1
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4029_ MuI._0339_ MuI._0570_ MuI._2975_ MuI._2976_ vssd1 vssd1 vccd1 vccd1 MuI._3129_
+ sky130_fd_sc_hd__nand4_1
XANTENNA__08134__C _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10680__B _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09825_ _02475_ _02476_ _02468_ _02473_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__o211ai_1
XANTENNA_input4_A Operation[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09756_ _02380_ _02387_ _02389_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__and3_1
X_06968_ _05080_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[17\] sky130_fd_sc_hd__buf_2
XANTENNA__06886__A _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08707_ _00950_ _01324_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__nor2_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _02153_ _02157_ _02327_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__and3_1
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _04338_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[6\] sky130_fd_sc_hd__clkbuf_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _01253_ _01255_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__or2_1
XFILLER_203_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4417__A2 MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11016__B _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07213__C _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ _01179_ _01180_ _01184_ _01185_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__or4_2
XFILLER_168_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ _03134_ _03298_ _03299_ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a31o_1
XFILLER_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07258__A2 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A1 _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _02712_ _03444_ _05948_ _06682_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__a22oi_1
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08455__B2 _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10262__A1 _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10531_ _03221_ _03236_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__nand3_1
XFILLER_183_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _02835_ _06095_ _02836_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__o21bai_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ _02987_ _04456_ _03160_ _03161_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__nand4_2
X_12201_ _04942_ _04808_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__a211o_1
XANTENNA__08758__A2 _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _05467_ _02945_ _06085_ _06086_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__a2111o_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10871__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _03085_ _03086_ _03088_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__and3_1
XFILLER_191_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12132_ _03378_ _00289_ _05252_ _05316_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__nand4_2
XFILLER_151_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1510_ AuI.pe.Significand\[0\] AuI._0695_ vssd1 vssd1 vccd1 vccd1 AuI._0696_
+ sky130_fd_sc_hd__or2_1
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ FuI.Integer\[12\] _02931_ _02938_ AuI.result\[12\] _04887_ vssd1 vssd1 vccd1
+ vccd1 _04888_ sky130_fd_sc_hd__a221o_1
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4709__B MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _00124_ _00125_ _06605_ _06591_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__and4_1
XAuI._1441_ AuI._0503_ AuI._0493_ vssd1 vssd1 vccd1 vccd1 AuI._0627_ sky130_fd_sc_hd__or2_1
XFILLER_93_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1372_ AuI._0389_ AuI._0471_ AuI._0422_ vssd1 vssd1 vccd1 vccd1 AuI._0564_ sky130_fd_sc_hd__and3_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06796__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0844__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ _05840_ _05841_ _05845_ _03315_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__a221o_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4380_ MuI._3342_ MuI._0061_ vssd1 vssd1 vccd1 vccd1 MuI._0062_ sky130_fd_sc_hd__xnor2_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _04724_ _04728_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand3_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _03346_ _05970_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__nand2_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _00877_ _00011_ _03444_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI._0860__A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6050_ MuI._1894_ MuI._1897_ vssd1 vssd1 vccd1 vccd1 MuI._1898_ sky130_fd_sc_hd__xnor2_1
XFILLER_199_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07249__A2 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._5001_ MuI._0741_ MuI._0742_ MuI._0743_ vssd1 vssd1 vccd1 vccd1 MuI._0744_ sky130_fd_sc_hd__o21bai_1
X_11778_ _04451_ _04453_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand2_1
XANTENNA__10253__A1 _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07420__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10253__B2 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729_ _02431_ _02229_ _03247_ _05820_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nand4_1
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08235__B _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13448_ _06358_ _06361_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__and2_1
XANTENNA__08749__A2 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ _06237_ _06241_ _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__o21a_1
XFILLER_142_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5903_ MuI._1698_ MuI._1700_ vssd1 vssd1 vccd1 vccd1 MuI._1737_ sky130_fd_sc_hd__and2b_1
XFILLER_154_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07421__A2 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5291__A MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5834_ MuI._1558_ MuI._1564_ MuI._1566_ vssd1 vssd1 vccd1 vccd1 MuI._1661_ sky130_fd_sc_hd__a21o_1
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09066__B _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _00041_ _00557_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__nor2_1
XFILLER_69_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._714_ AuI.pe._106_ AuI.pe._133_ AuI.pe._173_ AuI.pe._071_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._260_ sky130_fd_sc_hd__a22o_1
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5765_ MuI._2693_ MuI._2638_ MuI._2829_ MuI._3245_ vssd1 vssd1 vccd1 vccd1 MuI._1585_
+ sky130_fd_sc_hd__and4_1
XANTENNA__08401__D _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1639_ AuI.pe.Significand\[22\] AuI._0599_ AuI._0708_ AuI._0798_ AuI._0698_ vssd1
+ vssd1 vccd1 vccd1 AuI._0803_ sky130_fd_sc_hd__o221a_1
X_07871_ _00292_ _00301_ _00487_ _00488_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a22o_1
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6097__A1 MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6097__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._645_ AuI.pe._074_ AuI.pe._185_ AuI.pe._187_ AuI.pe._195_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[15\] sky130_fd_sc_hd__o22a_1
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4716_ MuI._1802_ MuI._0101_ MuI._3246_ MuI._2550_ vssd1 vssd1 vccd1 vccd1 MuI._0431_
+ sky130_fd_sc_hd__a22oi_1
X_09610_ _02205_ _00072_ _04434_ _06534_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
X_06822_ _03507_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__and3_1
XFILLER_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5696_ MuI._2873_ MuI._2785_ MuI._2875_ MuI._2765_ vssd1 vssd1 vccd1 vccd1 MuI._1509_
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._576_ AuI.pe._055_ AuI.pe._112_ AuI.pe._097_ AuI.pe._046_ AuI.pe._130_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._131_ sky130_fd_sc_hd__a221o_1
XFILLER_209_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4647_ MuI._0342_ MuI._0346_ MuI._0348_ vssd1 vssd1 vccd1 vccd1 MuI._0355_ sky130_fd_sc_hd__or3_1
X_09541_ _01332_ _02334_ _00592_ _00089_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__and4_1
XFILLER_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06753_ _02765_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__and3_1
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__B _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4578_ MuI._0270_ MuI._0271_ MuI._0278_ vssd1 vssd1 vccd1 vccd1 MuI._0279_ sky130_fd_sc_hd__a21bo_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _06488_ _04434_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nand2_1
XFILLER_24_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06684_ _02020_ net3 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__nor2_2
XMuI._6317_ MuI._2160_ MuI._2190_ vssd1 vssd1 vccd1 vccd1 MuI._2192_ sky130_fd_sc_hd__and2_1
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3529_ MuI._1164_ MuI._0526_ MuI._0757_ vssd1 vssd1 vccd1 vccd1 MuI._1175_ sky130_fd_sc_hd__and3_1
XANTENNA__09810__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ _00879_ _00876_ _00875_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5072__A2 MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6248_ MuI._0878_ MuI._3091_ MuI._2048_ MuI._2047_ vssd1 vssd1 vccd1 vccd1 MuI._2116_
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08354_ _00960_ _00959_ _00958_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__o21ai_1
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07305_ net40 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07330__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6179_ MuI._2023_ MuI._2032_ MuI._2031_ vssd1 vssd1 vccd1 vccd1 MuI._2040_ sky130_fd_sc_hd__a21o_1
XFILLER_165_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ _00900_ _00901_ _00891_ _00897_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__o211ai_2
XANTENNA_MuI._6021__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6021__B2 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ net130 vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__buf_4
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5780__B1 MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11787__A _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _06463_ _06461_ _05627_ _02107_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__a22oi_2
XFILLER_180_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__D _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07098_ _06412_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6297__A MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13497__A1 MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__B2 AuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12114__C _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _02418_ _02417_ _02416_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4099__B1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11953__C _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0972__A0 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07505__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _02309_ _02310_ _02311_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__or3_1
XFILLER_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _05622_ _05623_ _05613_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _04426_ _04427_ _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nand4_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _05549_ _05550_ _05512_ _05462_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__a211oi_1
XANTENNA_MuI._6260__A1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6260__B2 MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ _04383_ _04422_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or3_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08336__A _00951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__B1 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _02786_ _04326_ _01702_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o21a_1
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4711__C MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ _05724_ _02718_ _02731_ AuI.result\[26\] _06212_ vssd1 vssd1 vccd1 vccd1
+ _06213_ sky130_fd_sc_hd__a221o_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10514_ _03059_ _03061_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__nand2_1
XFILLER_183_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5095__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0941_ AuI._0152_ vssd1 vssd1 vccd1 vccd1 AuI._0153_ sky130_fd_sc_hd__buf_2
XFILLER_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _00345_ _04854_ _04274_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__a22o_1
XANTENNA__07651__A2 _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ _06139_ _06141_ _03133_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__o21ai_1
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__nor2_1
XAuI._0872_ AuI._0037_ AuI._0043_ AuI._0091_ vssd1 vssd1 vccd1 vccd1 AuI._0092_ sky130_fd_sc_hd__nand3_1
XFILLER_164_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10538__A2 _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0839__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08600__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13164_ _05751_ _05919_ _06064_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__o311a_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _02485_ _05638_ _06537_ _06565_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a22o_1
XMuI._3880_ MuI._2066_ MuI._2850_ MuI._2909_ MuI._2908_ vssd1 vssd1 vccd1 vccd1 MuI._2980_
+ sky130_fd_sc_hd__a31o_1
X_12115_ _03593_ _05025_ _06623_ net112 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__a22o_1
XFILLER_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13095_ _02782_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__or2_1
XANTENNA__10106__A _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._807__A AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12046_ _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__nand2_1
XFILLER_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07167__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07167__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5550_ MuI._1308_ MuI._1305_ MuI._1306_ vssd1 vssd1 vccd1 vccd1 MuI._1348_ sky130_fd_sc_hd__or3_1
XFILLER_77_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._526__B AuI.pe._070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1424_ AuI._0261_ AuI._0289_ AuI._0296_ AuI._0299_ vssd1 vssd1 vccd1 vccd1 AuI._0610_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12321__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._430_ AuI.pe._396_ vssd1 vssd1 vccd1 vccd1 AuI.pe._397_ sky130_fd_sc_hd__buf_2
XMuI._4501_ MuI._0078_ MuI._0193_ vssd1 vssd1 vccd1 vccd1 MuI._0194_ sky130_fd_sc_hd__xnor2_1
XMuI._5481_ MuI._1260_ MuI._1269_ MuI._1270_ MuI._1271_ vssd1 vssd1 vccd1 vccd1 MuI._1272_
+ sky130_fd_sc_hd__a211oi_4
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1355_ AuI._0547_ AuI._0548_ vssd1 vssd1 vccd1 vccd1 AuI._0549_ sky130_fd_sc_hd__nor2_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4432_ MuI._0094_ MuI._0095_ MuI._0117_ vssd1 vssd1 vccd1 vccd1 MuI._0118_ sky130_fd_sc_hd__nor3_1
XANTENNA__08116__B1 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1286_ AuI._0483_ AuI._0478_ vssd1 vssd1 vccd1 vccd1 AuI._0485_ sky130_fd_sc_hd__and2b_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _05835_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nand2_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4363_ MuI._3318_ MuI._3317_ vssd1 vssd1 vccd1 vccd1 MuI._0044_ sky130_fd_sc_hd__nor2_1
XFILLER_179_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _02805_ _05762_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__o21a_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5054__A2 MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6102_ MuI._1949_ MuI._1954_ vssd1 vssd1 vccd1 vccd1 MuI._1955_ sky130_fd_sc_hd__xnor2_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4294_ MuI._3310_ MuI._3311_ vssd1 vssd1 vccd1 vccd1 MuI._3394_ sky130_fd_sc_hd__and2_1
XFILLER_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13412__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6033_ MuI._1862_ MuI._1878_ vssd1 vssd1 vccd1 vccd1 MuI._1880_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4902__B MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12991__A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10777__A2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _00674_ _00675_ _00686_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__and3_1
XFILLER_140_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07021_ _05649_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11400__A _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08412__C _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6866_ MuI._2494_ MuI._0273_ vssd1 vssd1 vccd1 vccd1 MuI._2768_ sky130_fd_sc_hd__and2b_1
XFILLER_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _01566_ _01567_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__and4bb_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4349__B MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5817_ MuI._1556_ MuI._1641_ vssd1 vssd1 vccd1 vccd1 MuI._1642_ sky130_fd_sc_hd__xnor2_1
X_07923_ _06522_ _00535_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__nor2_1
XMuI._6797_ MuI._2685_ MuI._2596_ MuI._2600_ MuI._2697_ vssd1 vssd1 vccd1 vccd1 MuI._2720_
+ sky130_fd_sc_hd__or4_1
XFILLER_111_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5748_ MuI._1318_ MuI._1813_ MuI._0245_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._1566_
+ sky130_fd_sc_hd__and4_1
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07854_ _00455_ _00456_ _00471_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__nor3_1
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11773__C _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0889__A2_N net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._628_ AuI.pe._378_ AuI.pe._004_ AuI.pe._022_ AuI.pe._158_ AuI.pe._179_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._180_ sky130_fd_sc_hd__a221o_1
XANTENNA_AuI._0954__A0 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06805_ _03324_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__buf_4
XMuI._5679_ MuI._1487_ MuI._1488_ MuI._1489_ vssd1 vssd1 vccd1 vccd1 MuI._1490_ sky130_fd_sc_hd__nand3_1
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13046__B _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07785_ _00400_ _00401_ _00395_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a21o_1
XAuI.pe._559_ AuI.pe._030_ AuI.pe._112_ AuI.pe._079_ AuI.pe._046_ AuI.pe._115_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._116_ sky130_fd_sc_hd__a221o_1
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ _02149_ _02150_ _02152_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__nand3_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06736_ _02582_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__buf_6
XFILLER_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1596__A AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _02077_ _02078_ _06620_ _03873_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07979__B _00596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _02647_ _00032_ _06611_ _02582_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__a22o_1
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._110_ FuI._052_ FuI._056_ FuI.a_operand\[14\] vssd1 vssd1 vccd1 vccd1 FuI._004_
+ sky130_fd_sc_hd__o21a_1
X_09386_ _02002_ _02000_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08156__A _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08337_ _00817_ _00818_ _00954_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11414__B1 _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__C1 _05476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10768__A2 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ _00883_ _00884_ _00885_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__or3_1
XFILLER_165_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5346__D MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4250__D MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__buf_4
XFILLER_180_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08199_ _06458_ _00664_ _00663_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__nand3_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11310__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _02827_ _05724_ _02911_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o221a_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11193__A2 _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__A1 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _05531_ _03400_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and2b_1
XFILLER_161_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10940__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10092_ _02764_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__inv_2
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13237__A _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08897__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08897__B2 _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07235__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09153__C _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12802_ _03489_ _05672_ _05673_ _05676_ _05681_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__a311o_1
XAuI._1140_ AuI._0347_ AuI._0348_ vssd1 vssd1 vccd1 vccd1 AuI._0349_ sky130_fd_sc_hd__and2b_1
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ _03591_ _03594_ _03734_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__o211ai_1
XFILLER_71_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05605_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__xnor2_1
XAuI._1071_ net59 net27 net48 net16 AuI._0123_ AuI._0175_ vssd1 vssd1 vccd1 vccd1
+ AuI._0282_ sky130_fd_sc_hd__mux4_1
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _00292_ _03051_ _05530_ _05532_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__a22o_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3598__A2 MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11615_ _00132_ _00530_ _05445_ _00133_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a22oi_2
XANTENNA__11204__B _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _05440_ _05322_ _05458_ _05459_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a211o_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ FuI.Integer\[8\] _02931_ _02719_ _04542_ _04331_ vssd1 vssd1 vccd1 vccd1
+ _04332_ sky130_fd_sc_hd__a221o_1
XFILLER_156_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1673__A1 AuI._0116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10085__A_N _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0924_ AuI._0137_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[29\] sky130_fd_sc_hd__buf_2
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__B _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _06613_ _04255_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a21bo_1
XFILLER_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12316__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ _06122_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__and2_1
XMuI._4981_ MuI._0719_ MuI._0721_ vssd1 vssd1 vccd1 vccd1 MuI._0722_ sky130_fd_sc_hd__nand2_1
XFILLER_171_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _02752_ _02930_ _03127_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__a21o_2
XFILLER_125_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0855_ net11 net120 vssd1 vssd1 vccd1 vccd1 AuI._0075_ sky130_fd_sc_hd__and2b_1
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07388__A1 _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6720_ MuI._2241_ MuI._2634_ vssd1 vssd1 vccd1 vccd1 MuI._2635_ sky130_fd_sc_hd__xor2_1
XMuI._3932_ MuI._3020_ MuI._3024_ MuI._3018_ vssd1 vssd1 vccd1 vccd1 MuI._3032_ sky130_fd_sc_hd__o21a_1
XANTENNA__10481__D _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _05976_ _05978_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__and2b_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _02604_ _02669_ _06546_ _03051_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__nand4_1
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6651_ MuI._2513_ MuI._2542_ MuI._2544_ MuI._2558_ vssd1 vssd1 vccd1 vccd1 MuI._2559_
+ sky130_fd_sc_hd__or4_4
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3863_ MuI._2894_ MuI._2867_ MuI._2869_ MuI._0328_ vssd1 vssd1 vccd1 vccd1 MuI._2963_
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11874__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _05866_ _05880_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__or2_1
XMuI._5602_ MuI._1292_ MuI._1293_ MuI._1404_ vssd1 vssd1 vccd1 vccd1 MuI._1405_ sky130_fd_sc_hd__or3_1
XANTENNA_AuI._1189__A0 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12133__A1 _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3794_ MuI._0559_ vssd1 vssd1 vccd1 vccd1 MuI._2894_ sky130_fd_sc_hd__buf_2
XMuI._6582_ MuI._0691_ MuI._2478_ MuI._0548_ vssd1 vssd1 vccd1 vccd1 MuI._2483_ sky130_fd_sc_hd__a21oi_2
X_12029_ _04830_ _04849_ _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__and3_1
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0936__A0 net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5533_ MuI._1323_ MuI._1326_ MuI._1327_ MuI._1328_ vssd1 vssd1 vccd1 vccd1 MuI._1330_
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1407_ AuI._0594_ AuI._0595_ vssd1 vssd1 vccd1 vccd1 AuI._0596_ sky130_fd_sc_hd__or2_1
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._413_ AuI.pe.significand\[10\] vssd1 vssd1 vccd1 vccd1 AuI.pe._380_ sky130_fd_sc_hd__buf_2
XFILLER_53_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5464_ MuI._0100_ MuI._3262_ MuI._3397_ MuI._3362_ vssd1 vssd1 vccd1 vccd1 MuI._1254_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1338_ AuI._0482_ AuI._0530_ AuI._0531_ AuI._0533_ vssd1 vssd1 vccd1 vccd1 AuI._0534_
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _06661_ _06671_ _06670_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__a21o_1
XFILLER_207_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06984__A _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4415_ MuI.a_operand\[5\] vssd1 vssd1 vccd1 vccd1 MuI._0100_ sky130_fd_sc_hd__buf_2
XFILLER_207_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5395_ MuI._1176_ MuI._1177_ vssd1 vssd1 vccd1 vccd1 MuI._1178_ sky130_fd_sc_hd__xnor2_2
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1269_ AuI._0468_ AuI._0469_ vssd1 vssd1 vccd1 vccd1 AuI._0470_ sky130_fd_sc_hd__nand2_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4346_ MuI._0570_ MuI._3269_ vssd1 vssd1 vccd1 vccd1 MuI._0025_ sky130_fd_sc_hd__nand2_1
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _01262_ _01264_ _01266_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__o21a_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4277_ MuI._3375_ MuI._3376_ vssd1 vssd1 vccd1 vccd1 MuI._3377_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3589__A2 MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3529__A MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ _01717_ _01785_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__nand3_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1113__A0 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6016_ MuI._3098_ MuI._3100_ vssd1 vssd1 vccd1 vccd1 MuI._1861_ sky130_fd_sc_hd__and2_1
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _00737_ _00738_ _00739_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__and3_1
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._664__A_N AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _00499_ _00500_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout112_A net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07004_ _05467_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__and3_1
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5463__B MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6849_ MuI._2718_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[17\] sky130_fd_sc_hd__nor2_1
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08955_ _01255_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__nor2_1
XFILLER_130_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4710__A1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07906_ _00255_ _00370_ _00522_ _00523_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._4710__B2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _01498_ _01503_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08879__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07055__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09540__A2 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _00452_ _00453_ _00454_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__and3_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12896__A _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07768_ _00162_ _00163_ _00385_ _00164_ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a22oi_1
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06894__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _02130_ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__xor2_1
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06719_ _02399_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[5\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _00308_ _00315_ _00316_ _00298_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__o211ai_4
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__or2b_1
XFILLER_158_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _02474_ _00592_ _00089_ _06564_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07221__C _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _04327_ _02442_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or2b_1
XANTENNA__12060__B1 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _05226_ _05227_ _05146_ _05147_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__a211o_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ _00676_ _00048_ _00040_ _00506_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__a22o_1
XFILLER_193_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _03820_ _04391_ _03877_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__a31o_1
XFILLER_153_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11166__A2 _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ _05882_ _05811_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a21oi_1
X_10213_ _02893_ _02844_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o21ai_1
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _00058_ _05327_ _03949_ _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a22o_1
XFILLER_133_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input42_A b_operand[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _02820_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_95_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07891__C _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12115__B2 net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ _02735_ _02747_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__nor2_1
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10677__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5257__A2 MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__B _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1123_ AuI._0176_ AuI._0307_ AuI._0236_ AuI._0198_ AuI._0233_ vssd1 vssd1 vccd1
+ vccd1 AuI._0332_ sky130_fd_sc_hd__a41o_1
XANTENNA_MuI._5829__A MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09611__C _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10977_ _00289_ _00033_ _06612_ _00290_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__a22o_1
XFILLER_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4200_ MuI._3287_ MuI._3289_ MuI._3299_ vssd1 vssd1 vccd1 vccd1 MuI._3300_ sky130_fd_sc_hd__o21ai_2
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5180_ MuI._2799_ MuI._2918_ MuI._0110_ MuI.a_operand\[1\] vssd1 vssd1 vccd1
+ vccd1 MuI._0941_ sky130_fd_sc_hd__and4_1
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4217__B1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12716_ AuI.result\[18\] _02732_ _05586_ _05589_ vssd1 vssd1 vccd1 vccd1 _05590_
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1054_ AuI._0192_ AuI._0264_ vssd1 vssd1 vccd1 vccd1 AuI._0265_ sky130_fd_sc_hd__and2_1
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07845__A2 _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4131_ MuI._2807_ MuI._2806_ MuI._2794_ vssd1 vssd1 vccd1 vccd1 MuI._3231_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ _05513_ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__nor2_1
XFILLER_169_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08791__A2_N _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07131__C _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4062_ MuI._0350_ MuI._2967_ vssd1 vssd1 vccd1 vccd1 MuI._3162_ sky130_fd_sc_hd__nand2_1
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _05311_ _05317_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__nand2_1
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10601__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11529_ _04005_ _04153_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nor2_1
XFILLER_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0907_ net20 net114 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0127_ sky130_fd_sc_hd__mux2_1
XFILLER_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6098__C MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4964_ MuI._0618_ MuI._0703_ vssd1 vssd1 vccd1 vccd1 MuI._0704_ sky130_fd_sc_hd__nor2_1
XAuI._0838_ net116 net132 vssd1 vssd1 vccd1 vccd1 AuI._0058_ sky130_fd_sc_hd__or2b_1
XFILLER_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__A _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6703_ MuI._2604_ MuI._2615_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2617_ sky130_fd_sc_hd__mux2_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3915_ MuI._3013_ MuI._3014_ vssd1 vssd1 vccd1 vccd1 MuI._3015_ sky130_fd_sc_hd__nor2_1
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09355__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4895_ MuI._0619_ MuI._0627_ vssd1 vssd1 vccd1 vccd1 MuI._0628_ sky130_fd_sc_hd__xnor2_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6634_ MuI._2511_ MuI._2536_ MuI._2538_ MuI._2540_ vssd1 vssd1 vccd1 vccd1 MuI._2541_
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3846_ MuI._2385_ MuI._2407_ MuI._2396_ vssd1 vssd1 vccd1 vccd1 MuI._2946_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08740_ _01353_ _01357_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__xnor2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6565_ MuI._2461_ MuI._2463_ vssd1 vssd1 vccd1 vccd1 MuI._2465_ sky130_fd_sc_hd__and2_1
XMuI._3777_ MuI._1021_ MuI._2874_ MuI._2876_ MuI._0790_ vssd1 vssd1 vccd1 vccd1 MuI._2877_
+ sky130_fd_sc_hd__a22oi_1
X_08671_ _01285_ _01287_ _01288_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__a21bo_1
XFILLER_94_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5516_ MuI._1303_ MuI._1304_ MuI._1309_ vssd1 vssd1 vccd1 vccd1 MuI._1311_ sky130_fd_sc_hd__nand3_1
XFILLER_53_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07622_ _00236_ _00238_ _00239_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__nand3_1
XMuI._6496_ MuI._2243_ MuI._2305_ vssd1 vssd1 vccd1 vccd1 MuI._2389_ sky130_fd_sc_hd__or2_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08744__A2_N _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5447_ MuI._1229_ MuI._1233_ MuI._1234_ vssd1 vssd1 vccd1 vccd1 MuI._1235_ sky130_fd_sc_hd__o21ai_4
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07603__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0859__A1_N net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _00168_ _00169_ _00170_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__nand3_1
XFILLER_207_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4643__A MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5378_ MuI._1149_ MuI._1145_ vssd1 vssd1 vccd1 vccd1 MuI._1159_ sky130_fd_sc_hd__or2b_1
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07484_ _00092_ _00101_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4329_ MuI._3388_ MuI._0004_ MuI._0005_ vssd1 vssd1 vccd1 vccd1 MuI._0006_ sky130_fd_sc_hd__a21boi_1
X_09223_ _01758_ _01811_ _01840_ _01837_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a211o_1
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _01769_ _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10683__B _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11396__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ _00721_ _00719_ _00720_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__nand3_1
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09085_ _06516_ _00098_ _00047_ _06520_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a22oi_2
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08036_ _00652_ _00651_ _00650_ _00646_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__o211ai_2
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06889__A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09987_ _02651_ _02652_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08938_ _01554_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11019__B _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08869_ _06475_ _04907_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nand2_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _03632_ _03633_ _03460_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__a21bo_1
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ _04687_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__a21o_1
XFILLER_45_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07513__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _02948_ _06518_ _00412_ _02894_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a22o_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13073__A2 _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08884__A1_N _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5368__B MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ _03329_ _03485_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__nand2_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _05357_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__nor2_1
XFILLER_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10831__A1 _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _05992_ _02728_ _02931_ FuI.Integer\[31\] vssd1 vssd1 vccd1 vccd1 _06396_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10831__B2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _03410_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__nand3_2
XANTENNA__10874__A _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5411__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12432_ _05282_ _05283_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__and2b_1
XFILLER_139_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08899__A1_N _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08788__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _03733_ _05047_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__nand3_1
XFILLER_166_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09159__B _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10595__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08063__B _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11314_ _04078_ _04080_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__and3_1
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _05132_ _05135_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nand2_1
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12336__A1 _05092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11245_ _04005_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__or2_1
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1672_ AuI.exponent_sub\[7\] AuI._0695_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0023_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__06799__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10123__A_N _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10898__A1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _03786_ _03788_ _03787_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13409__B _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3700_ MuI._2799_ vssd1 vssd1 vccd1 vccd1 MuI._2800_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4728__A MuI.a_operand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08510__C _00896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4680_ MuI._0155_ MuI._0390_ vssd1 vssd1 vccd1 vccd1 MuI._0391_ sky130_fd_sc_hd__xnor2_1
X_10127_ _02801_ _05273_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__and2_1
XFILLER_110_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3631_ MuI._2209_ MuI._2275_ MuI._2286_ vssd1 vssd1 vccd1 vccd1 MuI._2297_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09504__A2 _01988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _02075_ _02729_ _02031_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__o21a_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6350_ MuI._2208_ MuI._2210_ MuI._2227_ vssd1 vssd1 vccd1 vccd1 MuI._2228_ sky130_fd_sc_hd__o21ba_1
XFILLER_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3562_ MuI._1340_ MuI._1527_ vssd1 vssd1 vccd1 vccd1 MuI._1538_ sky130_fd_sc_hd__nand2_1
XFILLER_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5301_ MuI._1070_ MuI._1072_ vssd1 vssd1 vccd1 vccd1 MuI._1074_ sky130_fd_sc_hd__xnor2_1
XMuI._3493_ MuI._0768_ vssd1 vssd1 vccd1 vccd1 MuI._0779_ sky130_fd_sc_hd__clkbuf_4
XMuI._6281_ MuI._2107_ MuI._2144_ vssd1 vssd1 vccd1 vccd1 MuI._2152_ sky130_fd_sc_hd__xor2_1
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5232_ MuI._0996_ MuI._0997_ vssd1 vssd1 vccd1 vccd1 MuI._0998_ sky130_fd_sc_hd__and2b_1
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1106_ AuI._0314_ AuI._0315_ AuI._0208_ vssd1 vssd1 vccd1 vccd1 AuI._0316_ sky130_fd_sc_hd__mux2_1
XANTENNA__12272__B1 _05092_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5163_ MuI._0919_ MuI._0920_ MuI._0912_ vssd1 vssd1 vccd1 vccd1 MuI._0923_ sky130_fd_sc_hd__a21o_1
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1037_ AuI._0110_ AuI._0248_ vssd1 vssd1 vccd1 vccd1 AuI._0249_ sky130_fd_sc_hd__xnor2_4
XFILLER_177_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4114_ MuI._2834_ MuI._3213_ vssd1 vssd1 vccd1 vccd1 MuI._3214_ sky130_fd_sc_hd__nand2_1
XMuI._5094_ MuI._0844_ MuI._0846_ vssd1 vssd1 vccd1 vccd1 MuI._0847_ sky130_fd_sc_hd__and2_1
XANTENNA__11599__B _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4045_ MuI._3142_ MuI._3143_ MuI._3144_ vssd1 vssd1 vccd1 vccd1 MuI._3145_ sky130_fd_sc_hd__nand3_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3807__A MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12207__C _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _02566_ _02568_ _02546_ _02569_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__and4bb_1
XMuI._5996_ MuI._0782_ MuI._1838_ vssd1 vssd1 vccd1 vccd1 MuI._1839_ sky130_fd_sc_hd__nor2_1
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4947_ MuI._0683_ MuI._0684_ MuI._2790_ MuI.b_operand\[8\] vssd1 vssd1 vccd1
+ vccd1 MuI._0685_ sky130_fd_sc_hd__and4bb_1
X_09841_ _02493_ _02494_ _02248_ _03960_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__and4bb_1
XFILLER_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4878_ MuI._0598_ MuI._0602_ MuI._0607_ MuI._0608_ vssd1 vssd1 vccd1 vccd1 MuI._0609_
+ sky130_fd_sc_hd__o211ai_2
X_09772_ _02414_ _02415_ _02419_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a21o_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _05252_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__clkbuf_4
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6617_ MuI._2521_ MuI._1452_ vssd1 vssd1 vccd1 vccd1 MuI._2522_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._3899__D MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3829_ MuI._1274_ MuI._2797_ vssd1 vssd1 vccd1 vccd1 MuI._2929_ sky130_fd_sc_hd__nand2_1
X_08723_ _01337_ _01340_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._731__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6548_ MuI._2438_ MuI._2441_ MuI._2439_ MuI._2432_ vssd1 vssd1 vccd1 vccd1 MuI._2446_
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08654_ _01245_ _01269_ _01271_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__o21a_1
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10678__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07605_ _00215_ _00220_ _00222_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__nand3_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6479_ MuI._1924_ MuI._1984_ MuI._2369_ vssd1 vssd1 vccd1 vccd1 MuI._2370_ sky130_fd_sc_hd__a21oi_1
X_08585_ _03239_ _03293_ _03884_ _03982_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__and4_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4373__A MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07536_ _06491_ net128 _00153_ _06492_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22oi_2
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4523__D MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10813__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ _00084_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__buf_4
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08482__A2 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _01693_ _01692_ _01685_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__a21o_1
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07398_ _00007_ _00008_ _00015_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nand3_1
XANTENNA__08164__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3717__A MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _01747_ _01750_ _01753_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a211oi_1
XANTENNA__10844__D _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0910__B_N net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10146__A_N _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5157__B2 MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _01596_ _01594_ _01595_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__or3_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08019_ _00540_ _00542_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10329__B1 _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08611__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _03772_ _03773_ _03617_ _03619_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o211a_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07508__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4548__A MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3452__A MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A2_N _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6185__D MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._722__A1 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12981_ _03497_ _05777_ _05871_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__and3_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10869__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11932_ _04744_ _04745_ _04589_ _04591_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o211ai_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07243__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11863_ _04670_ _04668_ _04669_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__nand3_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _02987_ _04596_ _03538_ _03540_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__nand4_2
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13451__C1 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11794_ _04554_ _04555_ _04595_ _04597_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10745_ _03243_ _03270_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13464_ _05992_ _02719_ _04642_ _05853_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a22o_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5826__B MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _03390_ _03391_ _03392_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a21o_1
XFILLER_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12308__B _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12415_ _05120_ _05122_ _05230_ _05231_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__o211a_1
XFILLER_173_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _05788_ _02726_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__nor2_1
XFILLER_182_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12346_ _05189_ _05190_ _05185_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21o_1
XANTENNA__08224__D _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__A _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0858__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__A1 _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5850_ MuI._1675_ MuI._1677_ vssd1 vssd1 vccd1 vccd1 MuI._1678_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12309__B2 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12277_ _05075_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__nand3_1
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._730_ AuI.pe._033_ AuI.pe._012_ AuI.pe._256_ AuI.pe._028_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._275_ sky130_fd_sc_hd__a22o_1
XMuI._4801_ MuI._0517_ MuI._0520_ MuI._0521_ MuI._0522_ vssd1 vssd1 vccd1 vccd1 MuI._0524_
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output73_A net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5781_ MuI._1600_ MuI._1601_ vssd1 vssd1 vccd1 vccd1 MuI._1602_ sky130_fd_sc_hd__nor2_1
X_11228_ _03812_ _03815_ _03987_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a211o_2
XANTENNA__07418__A _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1655_ AuI._0006_ AuI._0007_ AuI._0009_ vssd1 vssd1 vccd1 vccd1 AuI._0010_ sky130_fd_sc_hd__and3_1
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._661_ AuI.pe._196_ AuI.pe._198_ AuI.pe._207_ AuI.pe._210_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[16\] sky130_fd_sc_hd__o31a_1
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4732_ MuI._0878_ MuI._0246_ MuI._0446_ MuI._0447_ vssd1 vssd1 vccd1 vccd1 MuI._0448_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ _02442_ _05948_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__and3_1
XAuI._1586_ AuI._0259_ AuI._0758_ AuI._0759_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[11\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._592_ AuI.pe._145_ AuI.pe._141_ vssd1 vssd1 vccd1 vccd1 AuI.pe._146_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12978__B _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4663_ MuI._0246_ MuI._0471_ MuI._0239_ MuI._0242_ vssd1 vssd1 vccd1 vccd1 MuI._0373_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_AuI.pe._713__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6402_ MuI._2276_ MuI._2269_ MuI._2284_ vssd1 vssd1 vccd1 vccd1 MuI._2285_ sky130_fd_sc_hd__or3_1
XFILLER_209_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3614_ MuI._2011_ MuI._2099_ vssd1 vssd1 vccd1 vccd1 MuI._2110_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4594_ MuI._0219_ MuI._0290_ vssd1 vssd1 vccd1 vccd1 MuI._0297_ sky130_fd_sc_hd__nor2_1
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6333_ MuI._2169_ MuI._2183_ vssd1 vssd1 vccd1 vccd1 MuI._2210_ sky130_fd_sc_hd__nor2_1
XFILLER_36_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3545_ MuI._0592_ MuI._0889_ MuI._1197_ vssd1 vssd1 vccd1 vccd1 MuI._1351_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6264_ MuI._1043_ MuI._1285_ MuI._2016_ MuI._2014_ vssd1 vssd1 vccd1 vccd1 MuI._2134_
+ sky130_fd_sc_hd__a31o_1
XFILLER_211_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3476_ MuI._0581_ vssd1 vssd1 vccd1 vccd1 MuI._0592_ sky130_fd_sc_hd__buf_2
X_08370_ _06519_ net66 net11 net133 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__and4_1
XFILLER_205_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06992__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5215_ MuI._0842_ MuI._0979_ vssd1 vssd1 vccd1 vccd1 MuI._0980_ sky130_fd_sc_hd__or2_1
XFILLER_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ net38 vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__buf_4
XFILLER_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6195_ MuI._0361_ MuI._0603_ MuI._2849_ MuI._2914_ vssd1 vssd1 vccd1 vccd1 MuI._2058_
+ sky130_fd_sc_hd__and4_1
XANTENNA__08464__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5146_ MuI._0887_ MuI._0890_ MuI._0888_ vssd1 vssd1 vccd1 vccd1 MuI._0904_ sky130_fd_sc_hd__o21ba_1
XFILLER_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07252_ _06542_ _06543_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__nand3_1
XFILLER_177_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A1 _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5077_ MuI._0806_ MuI._0814_ MuI._0827_ vssd1 vssd1 vccd1 vccd1 MuI._0828_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07183_ _06478_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4028_ MuI._0790_ MuI._2851_ vssd1 vssd1 vccd1 vccd1 MuI._3128_ sky130_fd_sc_hd__nand2_1
XFILLER_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__D _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0815__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07328__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5979_ MuI._0771_ MuI._0772_ MuI._0774_ vssd1 vssd1 vccd1 vccd1 MuI._1820_ sky130_fd_sc_hd__a21o_1
XFILLER_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _02468_ _02473_ _02475_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a211o_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06967_ _05058_ _05069_ _04478_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__and3_1
X_09755_ _02391_ _02392_ _02387_ _02390_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__o211a_1
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08706_ _00947_ _00949_ _00948_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__o21a_1
X_09686_ _02153_ _02157_ _02327_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a21oi_1
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ _04327_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__and3_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _01253_ _01254_ _03002_ _00272_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__and4bb_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10201__B _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _01179_ _01180_ _01184_ _01185_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__o22ai_2
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07213__D _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__A1 _05559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07519_ _00094_ _00099_ _00097_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__o21bai_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08455__A2 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ _01116_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_211_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _03234_ _03235_ _03226_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a21o_1
XANTENNA__10262__A2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _02987_ _04456_ _03160_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a22o_1
XFILLER_136_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _03820_ _04865_ _04954_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__and3_1
X_13180_ _03400_ _05531_ _02721_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__o21a_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10392_ _03085_ _03086_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10871__B _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12131_ _00279_ _05252_ _00412_ _00278_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a22o_1
XFILLER_191_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09168__B1 _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ _04736_ _02727_ _02718_ _04800_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12711__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _01146_ _00550_ _00197_ _01147_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__a22oi_1
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4709__C MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1440_ AuI._0501_ AuI._0506_ vssd1 vssd1 vccd1 vccd1 AuI._0626_ sky130_fd_sc_hd__xnor2_2
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5302__A1 MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5302__B2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09453__A _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1371_ AuI._0556_ AuI._0563_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[19\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _02935_ _05847_ _05848_ _05850_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a311o_1
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _00345_ _05047_ _04726_ _04727_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__nand4_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12895_ _05692_ _05693_ _05733_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__nor3_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09900__B _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _04426_ _04498_ _04598_ _04599_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a211o_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04577_ _04578_ _04573_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4741__A MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5000_ MuI.a_operand\[17\] MuI.a_operand\[16\] MuI.b_operand\[1\] MuI.b_operand\[0\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0743_ sky130_fd_sc_hd__and4_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10253__A2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A1 _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _06560_ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__nand2_1
XANTENNA__07420__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13447_ _06358_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__nor2_1
X_10659_ _03355_ _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__xor2_2
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__nor2_1
XMuI._5902_ MuI._1733_ MuI._1734_ vssd1 vssd1 vccd1 vccd1 MuI._1735_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__or2_1
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5833_ MuI._1653_ MuI._1658_ vssd1 vssd1 vccd1 vccd1 MuI._1660_ sky130_fd_sc_hd__xnor2_2
XFILLER_170_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5291__B MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._713_ AuI.pe._056_ AuI.pe._089_ AuI.pe._197_ AuI.pe._150_ AuI.pe._102_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._259_ sky130_fd_sc_hd__a32o_1
XFILLER_123_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3552__B1 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5764_ MuI._2796_ MuI._0305_ vssd1 vssd1 vccd1 vccd1 MuI._1584_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._6330__A1_N MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1638_ AuI._0687_ AuI._0801_ AuI._0710_ vssd1 vssd1 vccd1 vccd1 AuI._0802_ sky130_fd_sc_hd__o21ai_1
X_07870_ _03378_ _00289_ _00074_ _00090_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__nand4_2
XAuI.pe._644_ AuI.pe._055_ AuI.pe._164_ AuI.pe._397_ AuI.pe._030_ AuI.pe._194_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._195_ sky130_fd_sc_hd__a221o_1
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4715_ MuI._3000_ MuI._2754_ MuI._2829_ MuI._0228_ vssd1 vssd1 vccd1 vccd1 MuI._0430_
+ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._6097__A2 MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06821_ _03497_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__clkbuf_4
XMuI._5695_ MuI._2790_ MuI._2867_ MuI._3223_ MuI._2875_ vssd1 vssd1 vccd1 vccd1 MuI._1508_
+ sky130_fd_sc_hd__nand4_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1569_ AuI._0639_ AuI._0745_ vssd1 vssd1 vccd1 vccd1 AuI._0746_ sky130_fd_sc_hd__xor2_1
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._575_ AuI.pe._028_ AuI.pe._119_ vssd1 vssd1 vccd1 vccd1 AuI.pe._130_ sky130_fd_sc_hd__and2_1
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4646_ MuI._0351_ MuI._0352_ MuI._0353_ vssd1 vssd1 vccd1 vccd1 MuI._0354_ sky130_fd_sc_hd__o21ba_1
X_09540_ _06504_ _04294_ _00072_ _06503_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06752_ _02754_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__buf_8
XFILLER_209_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13316__C _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4577_ MuI._0268_ MuI._0115_ MuI._0267_ vssd1 vssd1 vccd1 vccd1 MuI._0278_ sky130_fd_sc_hd__o21ai_1
X_09471_ _02092_ _02093_ _02091_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11117__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06683_ net4 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__buf_2
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6316_ MuI._2160_ MuI._2190_ vssd1 vssd1 vccd1 vccd1 MuI._2191_ sky130_fd_sc_hd__nor2_1
XFILLER_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3528_ MuI._1153_ vssd1 vssd1 vccd1 vccd1 MuI._1164_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ _00879_ _00875_ _00876_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__and3_1
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09810__B _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6247_ MuI._2113_ MuI._2114_ vssd1 vssd1 vccd1 vccd1 MuI._2115_ sky130_fd_sc_hd__nor2_1
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3459_ MuI.b_operand\[28\] MuI.b_operand\[27\] MuI.b_operand\[30\] MuI.b_operand\[29\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0405_ sky130_fd_sc_hd__or4_1
X_08353_ _00960_ _00958_ _00959_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__or3_1
XFILLER_211_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07304_ _06604_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__buf_4
XMuI._6178_ MuI._2035_ MuI._2038_ vssd1 vssd1 vccd1 vccd1 MuI._2039_ sky130_fd_sc_hd__or2b_1
XFILLER_177_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08284_ _00891_ _00897_ _00900_ _00901_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__a211o_1
XFILLER_177_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6021__A2 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5129_ MuI._0800_ MuI._0803_ MuI._0802_ vssd1 vssd1 vccd1 vccd1 MuI._0885_ sky130_fd_sc_hd__o21ba_1
XFILLER_137_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07235_ _02248_ _05638_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__nand2_1
XFILLER_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10972__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09538__A _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ _06460_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ _05134_ _06284_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._6297__B MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07058__A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4098__A MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13497__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06897__A _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09273__A _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _02418_ _02416_ _02417_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__or3_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4099__A1 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4099__B2 MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07999_ _03626_ _03928_ _04004_ _03561_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__a22o_4
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11953__D _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3730__A MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0972__A1 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _02376_ _02382_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__nor3_2
XANTENNA__10212__A _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__B1 _05160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__B _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ _02284_ _02286_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__xnor2_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11700_ _04291_ _04293_ _04475_ _04476_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__a211oi_2
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _05512_ _05462_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o211a_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08617__A _01233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6260__A2 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _04420_ _04421_ _04200_ _04384_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__o211a_1
XFILLER_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10484__A_N _03186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08336__B _00953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11562_ _02570_ _04347_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__nor2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _02705_ _02831_ _02832_ _02720_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a211oi_1
X_10513_ _03181_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__xor2_1
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4711__D MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0940_ AuI._0150_ AuI._0151_ vssd1 vssd1 vccd1 vccd1 AuI._0152_ sky130_fd_sc_hd__nand2_1
XFILLER_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _02983_ _02984_ _00550_ _04972_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__nand4_1
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13232_ _06063_ _06071_ _06061_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09448__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10444_ _06444_ _06442_ _00259_ _04369_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__and4_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0871_ AuI._0044_ net133 AuI._0045_ vssd1 vssd1 vccd1 vccd1 AuI._0091_ sky130_fd_sc_hd__o21ba_1
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _05915_ _05986_ _05987_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__o21ba_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ _05563_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__buf_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08600__A2 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ net112 _03593_ _05025_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__and3_1
XFILLER_124_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ _05994_ _02909_ _02926_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._4763__A1_N MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ _04864_ _04866_ _04867_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a21o_1
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07167__A2 _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0855__B net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1423_ AuI._0261_ AuI._0289_ AuI._0296_ AuI._0299_ vssd1 vssd1 vccd1 vccd1 AuI._0609_
+ sky130_fd_sc_hd__and4_1
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4500_ MuI._0080_ MuI._0079_ vssd1 vssd1 vccd1 vccd1 MuI._0193_ sky130_fd_sc_hd__nor2_1
XANTENNA__12321__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5480_ MuI._1202_ MuI._1213_ MuI._1212_ vssd1 vssd1 vccd1 vccd1 MuI._1271_ sky130_fd_sc_hd__a21oi_2
XFILLER_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1354_ AuI._0539_ AuI._0540_ AuI._0546_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0548_
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08116__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4431_ MuI._0115_ MuI._0116_ vssd1 vssd1 vccd1 vccd1 MuI._0117_ sky130_fd_sc_hd__or2_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1285_ AuI._0476_ AuI._0477_ vssd1 vssd1 vccd1 vccd1 AuI._0484_ sky130_fd_sc_hd__and2_1
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__inv_2
XFILLER_207_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4362_ MuI._0028_ MuI._0029_ MuI._0030_ vssd1 vssd1 vccd1 vccd1 MuI._0042_ sky130_fd_sc_hd__o21ba_1
XANTENNA_MuI._6787__A0 MuI._2563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13433__A _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6101_ MuI._1952_ MuI._1953_ vssd1 vssd1 vccd1 vccd1 MuI._1954_ sky130_fd_sc_hd__xnor2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _02805_ _05762_ _02711_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09383__A1_N _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4293_ MuI._3321_ MuI._3319_ vssd1 vssd1 vccd1 vccd1 MuI._3393_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11829_ _02926_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__buf_4
XANTENNA__13412__A2 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6032_ MuI._1872_ MuI._1877_ vssd1 vssd1 vccd1 vccd1 MuI._1878_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12991__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07020_ _05638_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__buf_4
XFILLER_162_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3815__A MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1443__A2 AuI._0519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6865_ MuI._2735_ MuI._2767_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[25\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__08412__D _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _01586_ _01587_ _01403_ _01413_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a211o_1
XMuI._5816_ MuI._1557_ MuI._1640_ vssd1 vssd1 vccd1 vccd1 MuI._1641_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6796_ MuI._2505_ MuI._2610_ MuI._2611_ vssd1 vssd1 vccd1 vccd1 MuI._2719_ sky130_fd_sc_hd__a21o_1
X_07922_ _00537_ _00539_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__nor2_1
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5747_ MuI._1558_ MuI._1564_ vssd1 vssd1 vccd1 vccd1 MuI._1565_ sky130_fd_sc_hd__xnor2_1
X_07853_ _00460_ _00470_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__xnor2_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI.pe._627_ AuI.pe._170_ AuI.pe._025_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._179_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__11773__D _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06804_ net114 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_AuI._0954__A1 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5678_ MuI._2851_ MuI._3247_ MuI._0997_ MuI._0996_ vssd1 vssd1 vccd1 vccd1 MuI._1489_
+ sky130_fd_sc_hd__a31o_1
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3828__A1 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _00395_ _00400_ _00401_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__and3_1
XANTENNA__12439__B1 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._558_ AuI.pe._084_ AuI.pe._042_ AuI.pe._097_ AuI.pe._013_ AuI.pe._114_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._115_ sky130_fd_sc_hd__a221o_1
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4629_ MuI._0332_ MuI._0334_ vssd1 vssd1 vccd1 vccd1 MuI._0335_ sky130_fd_sc_hd__or2b_1
XFILLER_83_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ _02149_ _02150_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a21o_1
X_06735_ net68 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07676__A2_N _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._540__C1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._489_ AuI.pe._020_ AuI.pe._050_ AuI.pe._042_ AuI.pe._029_ AuI.pe._051_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._052_ sky130_fd_sc_hd__a221o_1
XFILLER_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _06682_ _06436_ _06446_ _00000_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22oi_4
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08405_ _01019_ _01021_ _01020_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__o21ai_1
XANTENNA_MuI._4253__A1 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09385_ _02000_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__and2b_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08156__B _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08336_ _00951_ _00953_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__nand2_1
XANTENNA__11414__A1 _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5196__B MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__B1 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ _00062_ _04445_ _00085_ _00063_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__a22oi_1
XFILLER_119_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07218_ net107 vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__clkbuf_4
XFILLER_165_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09268__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08198_ _00814_ _00815_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__or2b_1
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11310__B _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _06429_ _03906_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__and3_1
XFILLER_134_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _03400_ _05531_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__and2b_1
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10091_ _02763_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__buf_2
XFILLER_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12422__A _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13237__B _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08897__A2 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__A _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07235__B _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09153__D _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12801_ _03110_ _02724_ _05677_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a211o_1
XFILLER_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _03731_ _03732_ _03713_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a21o_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ net114 _00385_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__and2_1
XAuI._1070_ AuI._0206_ AuI._0236_ AuI._0277_ AuI._0280_ vssd1 vssd1 vccd1 vccd1 AuI._0281_
+ sky130_fd_sc_hd__a31o_1
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _03486_ _05520_ _05530_ _05532_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nand4_1
XFILLER_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11614_ _04403_ _04404_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11204__C _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _05455_ _05457_ _05441_ _05442_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__o211a_1
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11545_ MuI.result\[8\] _02737_ _04011_ _04325_ _04330_ vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__a221o_1
XFILLER_184_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0923_ net26 net58 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0137_ sky130_fd_sc_hd__mux2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11476_ _03604_ _00033_ _06612_ _06434_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a22o_1
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12316__B _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3755__B1 MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4980_ MuI._0714_ MuI._0720_ vssd1 vssd1 vccd1 vccd1 MuI._0721_ sky130_fd_sc_hd__xnor2_1
X_10427_ _02933_ _02950_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or3_1
X_13215_ _03809_ _05660_ _06121_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a21o_1
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._0854_ net7 vssd1 vssd1 vccd1 vccd1 AuI._0074_ sky130_fd_sc_hd__inv_2
XFILLER_152_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3931_ MuI._3028_ MuI._3030_ vssd1 vssd1 vccd1 vccd1 MuI._3031_ sky130_fd_sc_hd__and2b_1
XANTENNA__07388__A2 _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _06682_ _06546_ _03051_ _00000_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a22o_1
X_13146_ _06047_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__xor2_1
XFILLER_152_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6650_ MuI._2551_ MuI._2557_ vssd1 vssd1 vccd1 vccd1 MuI._2558_ sky130_fd_sc_hd__or2_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3862_ MuI._0328_ MuI._2894_ MuI._2874_ MuI._2869_ vssd1 vssd1 vccd1 vccd1 MuI._2962_
+ sky130_fd_sc_hd__nand4_1
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13428__A _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__or2_1
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10289_ _00733_ _00741_ _00740_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a21o_1
XANTENNA__11874__C _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5601_ MuI._1333_ MuI._1403_ MuI._1330_ vssd1 vssd1 vccd1 vccd1 MuI._1404_ sky130_fd_sc_hd__a21o_1
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07139__A1_N _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1189__A1 net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12133__A2 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6581_ MuI._1747_ MuI._2308_ MuI._2475_ MuI._2477_ MuI._2481_ vssd1 vssd1 vccd1
+ vccd1 MuI._2482_ sky130_fd_sc_hd__o311a_2
X_12028_ _04847_ _04848_ _04735_ _04738_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a211o_1
XFILLER_211_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3793_ MuI._0328_ MuI._2892_ vssd1 vssd1 vccd1 vccd1 MuI._2893_ sky130_fd_sc_hd__and2_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4466__A MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5532_ MuI._1272_ MuI._1279_ MuI._1278_ vssd1 vssd1 vccd1 vccd1 MuI._1328_ sky130_fd_sc_hd__o21ai_1
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1406_ AuI.operand_a\[30\] AuI.exp_a AuI.operand_a\[24\] AuI.operand_a\[25\]
+ vssd1 vssd1 vccd1 vccd1 AuI._0595_ sky130_fd_sc_hd__or4_1
XANTENNA_AuI._0936__A1 net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._412_ AuI.pe._367_ AuI.pe._368_ AuI.pe._369_ AuI.pe._372_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._379_ sky130_fd_sc_hd__or4_2
XFILLER_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5463_ MuI._3268_ MuI._0228_ vssd1 vssd1 vccd1 vccd1 MuI._1253_ sky130_fd_sc_hd__nand2_1
XANTENNA__09641__A _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1337_ AuI._0521_ AuI._0532_ AuI._0529_ AuI._0511_ vssd1 vssd1 vccd1 vccd1 AuI._0533_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4414_ MuI.b_operand\[20\] MuI._3247_ vssd1 vssd1 vccd1 vccd1 MuI._0099_ sky130_fd_sc_hd__nand2_1
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5394_ MuI._1084_ MuI._1117_ MuI._1116_ vssd1 vssd1 vccd1 vccd1 MuI._1177_ sky130_fd_sc_hd__a21o_1
XAuI._1268_ AuI._0437_ AuI._0464_ AuI._0466_ AuI._0467_ vssd1 vssd1 vccd1 vccd1 AuI._0469_
+ sky130_fd_sc_hd__a31o_1
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08257__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__B2 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4345_ MuI._0019_ MuI._0023_ vssd1 vssd1 vccd1 vccd1 MuI._0024_ sky130_fd_sc_hd__or2_1
XANTENNA__07161__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1199_ AuI._0398_ AuI._0403_ AuI._0396_ vssd1 vssd1 vccd1 vccd1 AuI._0404_ sky130_fd_sc_hd__o21bai_2
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4276_ MuI._3367_ MuI._3374_ vssd1 vssd1 vccd1 vccd1 MuI._3376_ sky130_fd_sc_hd__or2_1
X_09170_ _02723_ _04186_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._3529__B MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__C _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6015_ MuI._1851_ MuI._1859_ vssd1 vssd1 vccd1 vccd1 MuI._1860_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1113__A1 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08121_ _00461_ _00463_ _00464_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__o21bai_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _00499_ _00500_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__nand2_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3746__B1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ _05456_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._5292__A2_N MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08720__A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__B1 _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6848_ MuI._2643_ MuI._2696_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[16\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_130_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08954_ _00058_ _00272_ _01253_ _01254_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4710__A2 MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6779_ MuI._2588_ MuI._2597_ MuI._2699_ MuI._2595_ vssd1 vssd1 vccd1 vccd1 MuI._2700_
+ sky130_fd_sc_hd__a22o_1
X_07905_ _00480_ _00481_ _00521_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__and3_1
XFILLER_97_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08885_ _01501_ _01502_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__nor2_1
XANTENNA__08879__A2 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07836_ _00214_ _00224_ _00223_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__a21bo_1
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12896__B _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._463__A AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07767_ net129 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _02131_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__xnor2_1
X_06718_ _02388_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__and3_1
XFILLER_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07839__B1 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08167__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07698_ _00265_ _00277_ _00297_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__or3_2
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09437_ _02046_ _02051_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__xnor2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__A1 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09368_ net106 _04229_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__and2_1
XFILLER_200_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07221__D _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12060__A1 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ _00891_ _00897_ _00900_ _00901_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a211oi_1
XFILLER_166_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _06631_ _06630_ _06436_ _06446_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__and4_1
XANTENNA__12417__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _00506_ _00676_ _00048_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__and3_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _03874_ _03876_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__nor2_1
XFILLER_180_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _02765_ _04736_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2b_1
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13000_ _05891_ _05892_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _00063_ _00062_ _05380_ _05445_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__nand4_1
XFILLER_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6151__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _03755_ _05917_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__nor2_1
XFILLER_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07891__D _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12115__A2 _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__A _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input35_A a_operand[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ MuI.result\[0\] _02739_ _06056_ FuI.Integer\[0\] _02746_ vssd1 vssd1 vccd1
+ vccd1 _02747_ sky130_fd_sc_hd__a221o_1
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._4717__C MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10677__A2 _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1122_ AuI._0180_ AuI._0185_ AuI._0187_ AuI._0292_ AuI._0206_ AuI._0189_ vssd1
+ vssd1 vccd1 vccd1 AuI._0331_ sky130_fd_sc_hd__mux4_1
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5829__B MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10976_ _03574_ _03577_ _03575_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21bai_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08077__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09611__D _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4217__A1 MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12715_ MuI.result\[18\] _02738_ _05587_ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_
+ sky130_fd_sc_hd__a211o_1
XAuI._1053_ AuI._0229_ AuI._0226_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0264_ sky130_fd_sc_hd__mux2_1
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4217__B2 MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4130_ MuI._2807_ MuI._2794_ MuI._2806_ vssd1 vssd1 vccd1 vccd1 MuI._3230_ sky130_fd_sc_hd__and3_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _06434_ _00678_ _00530_ _06666_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__and4_1
XFILLER_157_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07131__D _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08805__A _01419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4061_ MuI._2905_ MuI._2879_ MuI._2904_ vssd1 vssd1 vccd1 vccd1 MuI._3161_ sky130_fd_sc_hd__and3_1
XFILLER_169_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _05309_ _05171_ _05319_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__o21ai_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _04310_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__and2_1
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._0906_ AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0126_ sky130_fd_sc_hd__buf_4
X_11459_ _04230_ _04231_ _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or3b_1
XFILLER_125_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4963_ MuI._2583_ MuI._2830_ MuI._0616_ MuI._0617_ vssd1 vssd1 vccd1 vccd1 MuI._0703_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_MuI._6098__D MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0837_ net27 vssd1 vssd1 vccd1 vccd1 AuI._0057_ sky130_fd_sc_hd__inv_2
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08540__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3914_ MuI._2813_ MuI._2539_ MuI._2495_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._3014_
+ sky130_fd_sc_hd__a22oi_1
XMuI._6702_ MuI._2380_ MuI._2614_ vssd1 vssd1 vccd1 vccd1 MuI._2615_ sky130_fd_sc_hd__xor2_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4894_ MuI._0432_ MuI._0620_ vssd1 vssd1 vccd1 vccd1 MuI._0627_ sky130_fd_sc_hd__nor2_1
XANTENNA__09355__B _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13129_ _06029_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6633_ MuI._1712_ MuI._2537_ vssd1 vssd1 vccd1 vccd1 MuI._2540_ sky130_fd_sc_hd__nand2_1
XFILLER_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3845_ MuI._2943_ MuI._2944_ vssd1 vssd1 vccd1 vccd1 MuI._2945_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__A _06455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6564_ MuI._2461_ MuI._2463_ vssd1 vssd1 vccd1 vccd1 MuI._2464_ sky130_fd_sc_hd__nor2_1
XMuI._3776_ MuI._2875_ vssd1 vssd1 vccd1 vccd1 MuI._2876_ sky130_fd_sc_hd__buf_2
X_08670_ _01279_ _01284_ _01280_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI._1031__A0 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__A _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5515_ MuI._1303_ MuI._1304_ MuI._1309_ vssd1 vssd1 vccd1 vccd1 MuI._1310_ sky130_fd_sc_hd__a21o_1
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6495_ MuI._2307_ MuI._2337_ MuI._2387_ vssd1 vssd1 vccd1 vccd1 MuI._2388_ sky130_fd_sc_hd__or3_1
X_07621_ _03056_ _03099_ _00048_ _00033_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__nand4_1
XFILLER_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5446_ MuI._1161_ MuI._1168_ vssd1 vssd1 vccd1 vccd1 MuI._1234_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07552_ _00158_ _00159_ _00167_ vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4643__B MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5377_ MuI._1140_ MuI._1144_ vssd1 vssd1 vccd1 vccd1 MuI._1158_ sky130_fd_sc_hd__or2b_1
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07483_ _00094_ _00100_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4328_ MuI._0001_ MuI._0000_ MuI._0002_ vssd1 vssd1 vccd1 vccd1 MuI._0005_ sky130_fd_sc_hd__or3_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09222_ _01837_ _01809_ _01838_ _01839_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__nor4_2
XFILLER_210_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08715__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4259_ MuI._2817_ MuI._2330_ MuI._3237_ MuI._3238_ vssd1 vssd1 vccd1 vccd1 MuI._3359_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _02291_ _06548_ _00030_ _04703_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__and4_1
XFILLER_148_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08104_ _00719_ _00720_ _00721_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__a21o_1
XANTENNA__10683__C _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10053__B1 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _02528_ _00093_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nand2_4
XFILLER_175_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08035_ _00646_ _00650_ _00651_ _00652_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__a211o_2
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10980__A _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09986_ _01871_ _01213_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07066__A _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08937_ _01514_ _01516_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__nor2_1
XFILLER_130_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11019__C _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _01482_ _01484_ _01483_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a21o_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08721__A1 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09281__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__B2 _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07819_ _00408_ _00409_ _00435_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__nand3_1
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08799_ _06630_ _04176_ _04240_ _06631_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__a22oi_1
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _03419_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07513__B _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _03331_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5368__C MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _02703_ _04315_ _05356_ _04321_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a211oi_2
XANTENNA__10292__B1 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _06391_ _06393_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__nand2_2
X_10692_ _03393_ _03394_ _03410_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a21o_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__A2 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10874__B _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ _05279_ _05280_ _05281_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__a21o_1
XFILLER_166_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08788__A1 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5199__A2_N MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08788__B2 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12362_ _05207_ _05208_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10595__B2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__A _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _03967_ _03969_ _03968_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12293_ _05132_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__nor2_1
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11244_ _03657_ _03667_ _04006_ _03832_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__a31o_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1671_ AuI._0022_ vssd1 vssd1 vccd1 vccd1 AuI.result\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_122_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08360__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11544__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3913__A MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _03927_ _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10898__A2 _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0844__A_N net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _02801_ _05273_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__nor2_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10114__B _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3630_ MuI._2220_ MuI._2264_ vssd1 vssd1 vccd1 vccd1 MuI._2286_ sky130_fd_sc_hd__and2_1
X_10057_ net2 net1 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__and2_1
XFILLER_94_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3561_ MuI._1417_ MuI._1516_ vssd1 vssd1 vccd1 vccd1 MuI._1527_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07704__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5300_ MuI._1070_ MuI._1072_ vssd1 vssd1 vccd1 vccd1 MuI._1073_ sky130_fd_sc_hd__and2_1
XMuI._6280_ MuI._2149_ MuI._2150_ vssd1 vssd1 vccd1 vccd1 MuI._2151_ sky130_fd_sc_hd__xor2_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3492_ MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 MuI._0768_ sky130_fd_sc_hd__buf_2
XFILLER_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5231_ MuI._2837_ MuI.a_operand\[6\] MuI.a_operand\[5\] MuI.b_operand\[10\] vssd1
+ vssd1 vccd1 vccd1 MuI._0997_ sky130_fd_sc_hd__a22o_1
XANTENNA_AuI._1397__D AuI._0586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1105_ AuI._0230_ AuI._0239_ AuI._0223_ vssd1 vssd1 vccd1 vccd1 AuI._0315_ sky130_fd_sc_hd__mux2_1
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10959_ _03539_ _00678_ _00085_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__and3_1
XFILLER_16_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5162_ MuI._0912_ MuI._0919_ MuI._0920_ vssd1 vssd1 vccd1 vccd1 MuI._0921_ sky130_fd_sc_hd__nand3_1
XFILLER_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._550__B AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1036_ AuI._0157_ AuI._0159_ vssd1 vssd1 vccd1 vccd1 AuI._0248_ sky130_fd_sc_hd__and2_2
XFILLER_204_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6060__B1 MuI._1908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4113_ MuI._2809_ MuI._2810_ MuI._2833_ vssd1 vssd1 vccd1 vccd1 MuI._3213_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10784__B _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5093_ MuI._0795_ MuI._0843_ vssd1 vssd1 vccd1 vccd1 MuI._0846_ sky130_fd_sc_hd__nand2_1
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12629_ _00262_ _05895_ _05959_ _03110_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a22o_1
XANTENNA__11599__C _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4044_ MuI._3046_ MuI._3087_ vssd1 vssd1 vccd1 vccd1 MuI._3144_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._6603__A_N MuI._1836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3807__B MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11597__B1_N _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5995_ MuI._0673_ MuI._0781_ vssd1 vssd1 vccd1 vccd1 MuI._1838_ sky130_fd_sc_hd__and2_1
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4946_ MuI._0477_ MuI._3189_ MuI._3190_ MuI._0327_ vssd1 vssd1 vccd1 vccd1 MuI._0684_
+ sky130_fd_sc_hd__a22oi_1
X_09840_ _02205_ _06430_ _06431_ _06534_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a22oi_2
XANTENNA_AuI._1252__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4877_ MuI._0580_ MuI._0604_ MuI._0606_ vssd1 vssd1 vccd1 vccd1 MuI._0608_ sky130_fd_sc_hd__nand3_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09771_ _02416_ _02417_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__o21bai_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _05241_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__buf_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6616_ MuI._1453_ MuI._1372_ vssd1 vssd1 vccd1 vccd1 MuI._2521_ sky130_fd_sc_hd__or2b_1
XMuI._3828_ MuI._2860_ MuI._2914_ MuI._2920_ MuI._2917_ vssd1 vssd1 vccd1 vccd1 MuI._2928_
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08722_ _01338_ _01339_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__and2b_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1004__A0 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__A1 _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6547_ MuI._2424_ MuI._2444_ vssd1 vssd1 vccd1 vccd1 MuI._2445_ sky130_fd_sc_hd__nor2_1
XFILLER_67_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3759_ MuI._2847_ MuI._2848_ MuI._2857_ vssd1 vssd1 vccd1 vccd1 MuI._2859_ sky130_fd_sc_hd__a21o_1
X_08653_ _01157_ _01270_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10678__C _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6478_ MuI._1983_ MuI._1981_ vssd1 vssd1 vccd1 vccd1 MuI._2369_ sky130_fd_sc_hd__and2b_1
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _00221_ _06613_ _00218_ _00219_ vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__a22o_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _01188_ _01190_ _01191_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._4373__B MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5429_ MuI._1139_ MuI._1150_ MuI._1151_ vssd1 vssd1 vccd1 vccd1 MuI._1215_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI.pe._495__B2 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07535_ net28 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08467__B1 _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10274__B1 _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ net36 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__buf_2
XANTENNA__10813__A2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07987__C _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _01814_ _01821_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _00009_ _00014_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__xor2_1
XFILLER_195_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08164__B _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ _01434_ _01752_ _01729_ _01751_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__a211oi_1
XFILLER_194_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5157__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _01683_ _01684_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08018_ _00622_ _00634_ _00633_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__a21o_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10329__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08611__C _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07508__B _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09969_ _01676_ _01845_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__or2_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12980_ _03497_ _05777_ _05871_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__a21oi_1
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10869__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11931_ _04589_ _04591_ _04744_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a211o_1
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _04668_ _04669_ _04670_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__a21o_1
XFILLER_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._131__137 vssd1 vssd1 vccd1 vccd1 FuI._131__137/HI net137 sky130_fd_sc_hd__conb_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _03486_ _04596_ _03538_ _03540_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__a22o_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04554_ _04555_ _04595_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and4bb_1
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13261__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _03266_ _03269_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__nor2_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08355__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13463_ FuI.Integer\[30\] _02931_ _02938_ AuI.result\[30\] _06378_ vssd1 vssd1 vccd1
+ vccd1 _06379_ sky130_fd_sc_hd__a221o_1
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _03390_ _03391_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nand3_2
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12414_ _02865_ _05263_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__or2_1
XFILLER_154_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ _02707_ _02816_ _06307_ _02717_ _05853_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a32o_1
XANTENNA__10109__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _05185_ _05189_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nand3_2
XFILLER_127_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12309__A2 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08802__B _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12276_ _05114_ _05115_ _04975_ _05076_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__o211ai_1
XMuI._4800_ MuI._0517_ MuI._0520_ MuI._0521_ MuI._0522_ vssd1 vssd1 vccd1 vccd1 MuI._0523_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_135_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5780_ MuI._2765_ MuI._3189_ MuI._2875_ MuI._0477_ vssd1 vssd1 vccd1 vccd1 MuI._1601_
+ sky130_fd_sc_hd__a22oi_1
XAuI._1654_ AuI._0008_ AuI._0710_ vssd1 vssd1 vccd1 vccd1 AuI._0009_ sky130_fd_sc_hd__nand2_1
X_11227_ _03945_ _03946_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__o22a_1
XANTENNA__10125__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._660_ AuI.pe._208_ AuI.pe._209_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._210_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._6648__A2 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4731_ MuI._2939_ MuI._1142_ MuI._0305_ MuI._0445_ vssd1 vssd1 vccd1 vccd1 MuI._0447_
+ sky130_fd_sc_hd__and4_1
XANTENNA__12190__B1 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1585_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0760_ sky130_fd_sc_hd__buf_2
X_11158_ _02229_ _05884_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__and2_1
XANTENNA__07137__C net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._591_ AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 AuI.pe._145_ sky130_fd_sc_hd__buf_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4662_ MuI._0369_ MuI._0370_ vssd1 vssd1 vccd1 vccd1 MuI._0371_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ _02550_ _04467_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__and2b_1
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11089_ _02760_ _03838_ _02711_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6401_ MuI._2100_ MuI._2270_ vssd1 vssd1 vccd1 vccd1 MuI._2284_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI.pe._713__A2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3613_ MuI._2044_ MuI._2088_ vssd1 vssd1 vccd1 vccd1 MuI._2099_ sky130_fd_sc_hd__xor2_1
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4593_ MuI._0292_ MuI._0294_ vssd1 vssd1 vccd1 vccd1 MuI._0296_ sky130_fd_sc_hd__or2_1
XFILLER_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6332_ MuI._2168_ MuI._2167_ vssd1 vssd1 vccd1 vccd1 MuI._2208_ sky130_fd_sc_hd__and2b_1
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3544_ MuI._1285_ MuI._0526_ MuI._1329_ vssd1 vssd1 vccd1 vccd1 MuI._1340_ sky130_fd_sc_hd__and3_1
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6263_ MuI._2131_ MuI._2104_ vssd1 vssd1 vccd1 vccd1 MuI._2133_ sky130_fd_sc_hd__xnor2_1
XMuI._3475_ MuI._0570_ vssd1 vssd1 vccd1 vccd1 MuI._0581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__B2 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5214_ MuI._0828_ MuI._0841_ MuI._0837_ MuI._0840_ vssd1 vssd1 vccd1 vccd1 MuI._0979_
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13171__A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ _06620_ _05047_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__nand2_1
XFILLER_205_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6194_ MuI._0614_ MuI._2849_ MuI._2914_ MuI._0361_ vssd1 vssd1 vccd1 vccd1 MuI._2057_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_189_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5145_ MuI._0896_ MuI._0902_ vssd1 vssd1 vccd1 vccd1 MuI._0903_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07251_ _06547_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__xnor2_1
XAuI._1019_ AuI._0205_ AuI._0190_ AuI._0191_ AuI._0230_ vssd1 vssd1 vccd1 vccd1 AuI._0231_
+ sky130_fd_sc_hd__or4b_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5076_ MuI._0824_ MuI._0826_ vssd1 vssd1 vccd1 vccd1 MuI._0827_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__C _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07182_ _06481_ _06482_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__and2b_1
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4027_ MuI._3040_ MuI._3042_ MuI._3041_ vssd1 vssd1 vccd1 vccd1 MuI._3127_ sky130_fd_sc_hd__o21bai_1
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11756__B1 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09096__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__B1 _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5978_ MuI._1798_ MuI._1803_ MuI._1801_ vssd1 vssd1 vccd1 vccd1 MuI._1819_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07328__B _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4929_ MuI._0539_ MuI._0540_ vssd1 vssd1 vccd1 vccd1 MuI._0665_ sky130_fd_sc_hd__xor2_1
X_09823_ _02424_ _02433_ _02432_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._455__B AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._789_ AuI.pe._328_ AuI.pe._329_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[1\]
+ sky130_fd_sc_hd__nor2_1
X_09754_ _02401_ _02397_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__xor2_1
X_06966_ _02031_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__clkbuf_2
XFILLER_100_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08705_ _01196_ _01199_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__nand2_2
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _01919_ _02326_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__or2_1
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06897_ _04316_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__clkbuf_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08636_ _00062_ _04240_ _04305_ _00063_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__a22oi_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._468__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _01182_ _01183_ _01153_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__o21a_1
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10247__B1 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ _00130_ _00134_ _00131_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08498_ _01092_ _01105_ _01114_ _01115_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__a211oi_1
XFILLER_195_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07449_ _00057_ _00066_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _03389_ _02984_ _04520_ _00036_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand4_2
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._640__A1 AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _01427_ _01428_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10391_ _02259_ _05948_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__and3_1
XANTENNA__08612__B1 _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12425__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12130_ _04786_ _04788_ _04787_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__o21bai_1
XFILLER_151_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09168__A1 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3463__A MuI._0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09168__B2 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _00566_ _02745_ _04642_ _04671_ _04885_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a221o_1
XANTENNA__12172__B1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ _03751_ _03752_ _03753_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a21o_1
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4709__D MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1370_ AuI._0561_ AuI._0562_ vssd1 vssd1 vccd1 vccd1 AuI._0563_ sky130_fd_sc_hd__and2_1
XFILLER_65_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09453__B _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _05402_ _02719_ _05851_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a211o_1
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _03486_ _05047_ _04726_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a22o_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12894_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._812__C AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ _03831_ _04671_ _04568_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__nand3_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10131__B_N _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _04573_ _04577_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nand3_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4741__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ _06537_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11450__A2 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07420__C _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13446_ _06299_ _06360_ _06329_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21boi_1
X_10658_ _03372_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__nand2_1
XFILLER_139_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08603__B1 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _06275_ _06288_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and2_1
XFILLER_170_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _02562_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nor2_1
XMuI._5901_ MuI._1731_ MuI._1732_ MuI._1718_ MuI._1719_ vssd1 vssd1 vccd1 vccd1 MuI._1734_
+ sky130_fd_sc_hd__a211o_1
XFILLER_127_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07429__A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ _05163_ _05170_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__nor2_1
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10961__A1 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5832_ MuI._1654_ MuI._1657_ vssd1 vssd1 vccd1 vccd1 MuI._1658_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5291__C MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12259_ _02987_ _05262_ _05095_ _05096_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nand4_1
XFILLER_123_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._712_ AuI.pe._084_ AuI.pe._164_ AuI.pe._225_ AuI.pe._055_ AuI.pe._257_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._258_ sky130_fd_sc_hd__a221o_1
XANTENNA_MuI._3552__A1 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5763_ MuI._1578_ MuI._1579_ MuI._1580_ vssd1 vssd1 vccd1 vccd1 MuI._1583_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1637_ AuI._0686_ AuI._0690_ AuI._0688_ vssd1 vssd1 vccd1 vccd1 AuI._0801_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._643_ AuI.pe._063_ AuI.pe._119_ AuI.pe._188_ AuI.pe._193_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._194_ sky130_fd_sc_hd__a211o_1
XMuI._4714_ MuI._0294_ MuI._0426_ MuI._0428_ vssd1 vssd1 vccd1 vccd1 MuI._0429_ sky130_fd_sc_hd__or3_1
XMuI._5694_ MuI._0168_ MuI._3349_ vssd1 vssd1 vccd1 vccd1 MuI._1507_ sky130_fd_sc_hd__nand2_1
X_06820_ _03486_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1568_ AuI._0635_ AuI._0636_ AuI._0736_ AuI._0637_ vssd1 vssd1 vccd1 vccd1 AuI._0745_
+ sky130_fd_sc_hd__o31a_1
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4645_ MuI.a_operand\[15\] MuI.a_operand\[14\] MuI._2866_ MuI.b_operand\[6\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0353_ sky130_fd_sc_hd__and4_1
XAuI.pe._574_ AuI.pe._122_ AuI.pe._124_ AuI.pe._128_ AuI.pe._129_ AuI.pe._074_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe.Significand\[10\] sky130_fd_sc_hd__o32a_1
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06751_ net40 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__buf_4
XAuI._1499_ AuI._0680_ AuI._0682_ vssd1 vssd1 vccd1 vccd1 AuI._0685_ sky130_fd_sc_hd__nand2_1
XFILLER_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13316__D _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4576_ MuI._0275_ MuI._0276_ vssd1 vssd1 vccd1 vccd1 MuI._0277_ sky130_fd_sc_hd__xnor2_1
X_09470_ _02091_ _02092_ _02093_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__or3_1
XFILLER_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3527_ MuI._1142_ vssd1 vssd1 vccd1 vccd1 MuI._1153_ sky130_fd_sc_hd__buf_2
XMuI._6315_ MuI._2188_ MuI._2189_ vssd1 vssd1 vccd1 vccd1 MuI._2190_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ _00855_ _01036_ _01037_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__a21o_1
XFILLER_197_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09810__C net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6246_ MuI._0878_ MuI._2077_ MuI._2112_ vssd1 vssd1 vccd1 vccd1 MuI._2114_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3458_ MuI._0350_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._0394_ sky130_fd_sc_hd__and2_1
X_08352_ _00963_ _00964_ _00969_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__nand3_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6177_ MuI._2035_ MuI._2036_ MuI._2037_ vssd1 vssd1 vccd1 vccd1 MuI._2038_ sky130_fd_sc_hd__or3_1
X_07303_ net11 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ _00899_ _00898_ _00868_ _00866_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__o211a_1
XFILLER_192_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5128_ MuI._0881_ MuI._0882_ MuI._0865_ vssd1 vssd1 vccd1 vccd1 MuI._0884_ sky130_fd_sc_hd__a21o_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07234_ _06534_ _06491_ net130 net129 vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__and4_1
XFILLER_165_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10972__B _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1374__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5059_ MuI._2873_ MuI._3190_ MuI.a_operand\[5\] MuI._3245_ vssd1 vssd1 vccd1
+ vccd1 MuI._0808_ sky130_fd_sc_hd__nand4_1
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ net21 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._5780__A2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__B _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3791__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12941__A2 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _06411_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6297__C MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4098__B MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09806_ _02456_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__nor2_1
XFILLER_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09273__B _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4099__A2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07998_ _00317_ _00613_ _00612_ _00602_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__a211o_1
XANTENNA__07581__B1 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07074__A _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09737_ _02307_ _02375_ _02366_ _02374_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a211oi_2
XANTENNA__12457__A1 _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _04876_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[14\] sky130_fd_sc_hd__clkbuf_2
X_09668_ _02304_ _02307_ _02256_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a211oi_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _01235_ _01232_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09599_ _02168_ _02169_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _04200_ _04384_ _04420_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__a211oi_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3458__A MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11561_ _02546_ _02548_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11432__A2 _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ MuI.result\[26\] _02738_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a21o_1
XFILLER_195_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _03215_ _03216_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__nand2_1
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5220__A1 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11492_ _02980_ _04907_ _04972_ _00281_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5673__A MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13231_ _06137_ _06138_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__or2b_1
XFILLER_183_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10443_ _03615_ _00259_ _04369_ _03550_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__a22oi_1
XAuI._0870_ AuI._0077_ AuI._0088_ AuI._0089_ AuI._0075_ vssd1 vssd1 vccd1 vccd1 AuI._0090_
+ sky130_fd_sc_hd__o22a_1
XFILLER_183_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input65_A b_operand[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _05918_ _05988_ _05921_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or3b_1
X_10374_ _00782_ _00784_ _00786_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o21bai_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10943__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ _04770_ _04804_ _04805_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or3_1
XFILLER_124_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13093_ _02908_ _05859_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12044_ _04864_ _04866_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nand3_1
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1422_ AuI._0253_ AuI._0607_ vssd1 vssd1 vccd1 vccd1 AuI._0608_ sky130_fd_sc_hd__and2_1
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07572__B1 _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12321__C _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1353_ AuI._0539_ AuI._0540_ AuI._0546_ vssd1 vssd1 vccd1 vccd1 AuI._0547_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._137__143 vssd1 vssd1 vccd1 vccd1 FuI._137__143/HI net143 sky130_fd_sc_hd__conb_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6009__A MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4430_ MuI._0105_ MuI._0114_ vssd1 vssd1 vccd1 vccd1 MuI._0116_ sky130_fd_sc_hd__nor2_1
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08116__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B1 _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1284_ AuI._0478_ AuI._0483_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[12\]
+ sky130_fd_sc_hd__xnor2_4
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12946_ _05740_ _05776_ _05834_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__and3_1
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07324__B1 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4361_ MuI._0038_ MuI._0039_ MuI._0040_ vssd1 vssd1 vccd1 vccd1 MuI._0041_ sky130_fd_sc_hd__o21ba_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6100_ MuI._2791_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._1953_ sky130_fd_sc_hd__nand2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _05581_ _05759_ _05760_ _05761_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4292_ MuI._3338_ MuI._3391_ vssd1 vssd1 vccd1 vccd1 MuI._3392_ sky130_fd_sc_hd__and2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _02860_ _04493_ _02858_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6031_ MuI._1875_ MuI._1876_ vssd1 vssd1 vccd1 vccd1 MuI._1877_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1429__B_N AuI._0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12620__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__xor2_4
XFILLER_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09639__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__B _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13429_ _01320_ _06305_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nand2_1
XFILLER_127_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07159__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3815__B MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0999_ AuI._0096_ AuI._0150_ AuI._0156_ vssd1 vssd1 vccd1 vccd1 AuI._0211_ sky130_fd_sc_hd__nand3_1
XFILLER_170_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6864_ MuI._2766_ MuI._2491_ vssd1 vssd1 vccd1 vccd1 MuI._2767_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4870__A1_N MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _01403_ _01413_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__o211ai_2
XANTENNA__06998__A _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5815_ MuI._1638_ MuI._1639_ vssd1 vssd1 vccd1 vccd1 MuI._1640_ sky130_fd_sc_hd__nor2_1
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07921_ _00537_ _00538_ _06663_ _06584_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__and4bb_1
XMuI._6795_ MuI._2643_ MuI._2647_ vssd1 vssd1 vccd1 vccd1 MuI._2718_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5746_ MuI._1559_ MuI._1563_ vssd1 vssd1 vccd1 vccd1 MuI._1564_ sky130_fd_sc_hd__xnor2_2
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07852_ _00468_ _00469_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__and2b_1
XAuI.pe._626_ AuI.pe._089_ AuI.pe._086_ AuI.pe._053_ AuI.pe._125_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._178_ sky130_fd_sc_hd__a22o_1
XFILLER_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06803_ _03304_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[22\] sky130_fd_sc_hd__clkbuf_2
Xinput1 Operation[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XMuI._5677_ MuI._1485_ MuI._1486_ MuI._1484_ vssd1 vssd1 vccd1 vccd1 MuI._1488_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12439__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3828__A2 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07783_ _00397_ _00399_ _00396_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12439__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._557_ AuI.pe._071_ AuI.pe._004_ AuI.pe._023_ AuI.pe._393_ AuI.pe._113_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._114_ sky130_fd_sc_hd__a221o_1
XMuI._4628_ MuI._0184_ MuI._0333_ vssd1 vssd1 vccd1 vccd1 MuI._0334_ sky130_fd_sc_hd__xnor2_1
X_09522_ _02004_ _02007_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__xnor2_1
X_06734_ _02561_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[8\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_AuI.pe._540__B1 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4559_ MuI._0255_ MuI._0202_ MuI._0257_ vssd1 vssd1 vccd1 vccd1 MuI._0258_ sky130_fd_sc_hd__a21oi_1
XAuI.pe._488_ AuI.pe._033_ AuI.pe._023_ AuI.pe._027_ AuI.pe._045_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._051_ sky130_fd_sc_hd__a22o_1
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _02593_ _06583_ _06436_ _06430_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__and4_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08404_ _01019_ _01020_ _01021_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__or3_1
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09384_ _01901_ _02001_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__nor2_1
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6229_ MuI._2093_ MuI._2094_ vssd1 vssd1 vccd1 vccd1 MuI._2095_ sky130_fd_sc_hd__nor2_1
XANTENNA__08156__C _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08335_ _00661_ _00952_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__nor2_2
XANTENNA__08815__B1 _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5196__C MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1667__B1 AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ net119 _00090_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__nand2_1
XFILLER_192_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08453__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07217_ net17 vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__buf_6
XANTENNA__09268__B _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08197_ _00813_ _00665_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__or2b_1
XFILLER_180_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07148_ _06441_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__xor2_1
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09240__B1 _01266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ _06264_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10090_ _02761_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__or2_1
XANTENNA__06701__A _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4837__A MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__B _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3741__A MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A1 _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__B _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ FuI.Integer\[19\] _04627_ _02718_ _05273_ _05679_ vssd1 vssd1 vccd1 vccd1
+ _05680_ sky130_fd_sc_hd__a221o_1
XFILLER_28_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._531__B1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10992_ _03713_ _03731_ _03732_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nand3_1
XANTENNA__07306__B1 _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08628__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07532__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12731_ _05602_ _05603_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__o21ai_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11054__A _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ _03378_ _00289_ _03424_ _00382_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__nand4_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _00270_ _00423_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__nand2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12593_ _05441_ _05442_ _05455_ _05457_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__a211oi_4
XFILLER_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11204__D _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _02550_ _04467_ _02743_ _02944_ _04391_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a32o_1
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0814__C_N net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3916__A MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0922_ AuI._0136_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[28\] sky130_fd_sc_hd__clkbuf_2
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ _06434_ _03604_ _00033_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__and3_1
XFILLER_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3755__A1 MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3755__B2 MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._099_ FuI._037_ FuI._056_ FuI._058_ vssd1 vssd1 vccd1 vccd1 FuI._059_ sky130_fd_sc_hd__and3_1
XANTENNA__12316__C _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13214_ _03809_ _05671_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__nand3_1
X_10426_ _06428_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nor2_1
XFILLER_152_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0853_ AuI._0068_ net10 AuI._0071_ net9 vssd1 vssd1 vccd1 vccd1 AuI._0073_ sky130_fd_sc_hd__o22a_1
XANTENNA__10117__B _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3930_ MuI._2937_ MuI._2951_ MuI._3029_ vssd1 vssd1 vccd1 vccd1 MuI._3030_ sky130_fd_sc_hd__o21ai_2
XFILLER_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ _05940_ _06048_ _05974_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__a21o_1
XFILLER_112_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ _05498_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08810__B _01422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3861_ MuI._0779_ MuI._2871_ vssd1 vssd1 vccd1 vccd1 MuI._2961_ sky130_fd_sc_hd__nand2_1
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _05954_ _05973_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nor2_1
X_10288_ _02975_ _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__xnor2_4
XMuI._5600_ MuI._1365_ MuI._1367_ MuI._1368_ MuI._1369_ vssd1 vssd1 vccd1 vccd1 MuI._1403_
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11874__D _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1043__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3792_ MuI._2884_ vssd1 vssd1 vccd1 vccd1 MuI._2892_ sky130_fd_sc_hd__clkbuf_4
XMuI._6580_ MuI._2479_ MuI._2480_ vssd1 vssd1 vccd1 vccd1 MuI._2481_ sky130_fd_sc_hd__or2_1
XFILLER_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12027_ _04735_ _04738_ _04847_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o211ai_2
XANTENNA_MuI._4466__B MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5531_ MuI._1272_ MuI._1278_ MuI._1279_ vssd1 vssd1 vccd1 vccd1 MuI._1327_ sky130_fd_sc_hd__or3_1
XFILLER_66_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1405_ AuI.operand_a\[26\] AuI.operand_a\[27\] AuI.operand_a\[28\] AuI.operand_a\[29\]
+ vssd1 vssd1 vccd1 vccd1 AuI._0594_ sky130_fd_sc_hd__or4_1
XAuI.pe._411_ AuI.pe.significand\[11\] vssd1 vssd1 vccd1 vccd1 AuI.pe._378_ sky130_fd_sc_hd__buf_2
XFILLER_65_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5462_ MuI._1196_ MuI._1195_ MuI._1194_ vssd1 vssd1 vccd1 vccd1 MuI._1251_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09641__B _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1336_ AuI._0507_ AuI._0520_ vssd1 vssd1 vccd1 vccd1 AuI._0532_ sky130_fd_sc_hd__nor2_1
XANTENNA__07293__A1_N _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B1 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4413_ MuI._3361_ MuI._0096_ vssd1 vssd1 vccd1 vccd1 MuI._0098_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5393_ MuI._1173_ MuI._1174_ vssd1 vssd1 vccd1 vccd1 MuI._1176_ sky130_fd_sc_hd__nor2_1
XANTENNA__07442__A _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12929_ _05813_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1267_ AuI._0437_ AuI._0464_ AuI._0466_ AuI._0467_ vssd1 vssd1 vccd1 vccd1 AuI._0468_
+ sky130_fd_sc_hd__nand4_1
XFILLER_179_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11644__A2 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4344_ MuI._0019_ MuI._0022_ MuI._0768_ MuI._3268_ vssd1 vssd1 vccd1 vccd1 MuI._0023_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__12192__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08257__B _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07161__B _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1198_ AuI._0398_ AuI._0403_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[6\]
+ sky130_fd_sc_hd__xor2_2
XFILLER_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4275_ MuI._3367_ MuI._3374_ vssd1 vssd1 vccd1 vccd1 MuI._3375_ sky130_fd_sc_hd__nand2_1
XANTENNA__13397__A2 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6014_ MuI._1852_ MuI._1858_ vssd1 vssd1 vccd1 vccd1 MuI._1859_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08120_ _00734_ _00735_ _00736_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ _00482_ _00667_ _00668_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a21bo_2
XFILLER_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._3746__A1 MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ _05445_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08720__B _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__A1 _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6847_ MuI._2756_ vssd1 vssd1 vccd1 vccd1 MuI._2757_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__B2 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _01522_ _01524_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__nor2_1
XFILLER_102_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07904_ _00480_ _00481_ _00521_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__a21oi_2
XMuI._6778_ MuI._2685_ MuI._2591_ vssd1 vssd1 vccd1 vccd1 MuI._2699_ sky130_fd_sc_hd__or2_1
XANTENNA__10043__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _06663_ _00033_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07536__B1 _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__A1 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5729_ MuI._1052_ MuI._1479_ MuI._1543_ MuI._1544_ vssd1 vssd1 vccd1 vccd1 MuI._1545_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_111_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ _00450_ _00451_ _00442_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__a21o_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._609_ AuI.pe._072_ AuI.pe._086_ AuI.pe._157_ AuI.pe._161_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._162_ sky130_fd_sc_hd__a211o_1
XANTENNA__10978__A _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5120__B1 MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07766_ _06503_ _06504_ net130 net129 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__and4_1
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09505_ _01986_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06717_ _02377_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__buf_4
XANTENNA__07839__A1 _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07839__B2 _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07697_ _00313_ _00314_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__and2b_1
XFILLER_198_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09436_ _02054_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__nor2_1
XANTENNA__10843__B1 _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5423__A1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5423__B2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _01982_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _00934_ _00935_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__or2_1
XFILLER_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12060__A2 _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _00011_ _03960_ _06446_ _00012_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3736__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _00863_ _00864_ _00865_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__nand3_1
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0863__B2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ _04001_ _04003_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__or2_1
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10211_ _02878_ _02892_ _02870_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09726__B _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _00046_ _00530_ _06666_ _00049_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a22o_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11571__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _02818_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._6151__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3471__A MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _02741_ _02745_ _02559_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07246__B _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4717__D MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A a_operand[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10888__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1121_ AuI._0209_ vssd1 vssd1 vccd1 vccd1 AuI._0330_ sky130_fd_sc_hd__buf_2
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10975_ _03578_ _03586_ _03585_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__a21o_1
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08077__B _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12714_ FuI.Integer\[18\] _06045_ _02718_ _05209_ vssd1 vssd1 vccd1 vccd1 _05588_
+ sky130_fd_sc_hd__a22o_1
XAuI._1052_ AuI._0262_ vssd1 vssd1 vccd1 vccd1 AuI._0263_ sky130_fd_sc_hd__buf_2
XFILLER_31_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4217__A2 MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ _00676_ _05380_ _05445_ _00506_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a22oi_1
XFILLER_157_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6721__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4060_ MuI._3079_ MuI._3159_ vssd1 vssd1 vccd1 vccd1 MuI._3160_ sky130_fd_sc_hd__nand2_2
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12576_ _05437_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10062__A1 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11527_ _04307_ _04309_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand2_1
XFILLER_157_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output96_A net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0905_ AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0125_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ _04234_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0877__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08591__A1_N _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4962_ MuI._0699_ MuI._0697_ vssd1 vssd1 vccd1 vccd1 MuI._0701_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10409_ _03104_ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__xnor2_2
XFILLER_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0836_ AuI._0049_ AuI._0052_ AuI._0055_ vssd1 vssd1 vccd1 vccd1 AuI._0056_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11389_ _02771_ _02772_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__nand2_1
XMuI._6701_ MuI._2391_ MuI._2613_ vssd1 vssd1 vccd1 vccd1 MuI._2614_ sky130_fd_sc_hd__nor2_1
XANTENNA__08540__B _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3913_ MuI._2939_ MuI._2811_ MuI._2451_ MuI._2495_ vssd1 vssd1 vccd1 vccd1 MuI._3013_
+ sky130_fd_sc_hd__and4_1
XFILLER_152_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _05961_ _05964_ _06028_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand3_1
XMuI._4893_ MuI._0622_ MuI._0624_ vssd1 vssd1 vccd1 vccd1 MuI._0626_ sky130_fd_sc_hd__or2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4477__A MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6632_ MuI._1712_ MuI._2537_ vssd1 vssd1 vccd1 vccd1 MuI._2538_ sky130_fd_sc_hd__or2_1
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4908__C MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3844_ MuI._2812_ MuI._2816_ vssd1 vssd1 vccd1 vccd1 MuI._2944_ sky130_fd_sc_hd__nor2_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _03615_ _05713_ _05777_ _03550_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a22o_1
XANTENNA__07156__B _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3775_ MuI._2868_ vssd1 vssd1 vccd1 vccd1 MuI._2875_ sky130_fd_sc_hd__clkbuf_4
XMuI._6563_ MuI._2235_ MuI._2237_ vssd1 vssd1 vccd1 vccd1 MuI._2463_ sky130_fd_sc_hd__nor2_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1031__A1 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10798__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5514_ MuI._1305_ MuI._1306_ MuI._1308_ vssd1 vssd1 vccd1 vccd1 MuI._1309_ sky130_fd_sc_hd__o21bai_1
X_07620_ _00081_ _04638_ _04703_ _00237_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__a22o_1
XMuI._6494_ MuI._2338_ MuI._2364_ vssd1 vssd1 vccd1 vccd1 MuI._2387_ sky130_fd_sc_hd__nor2_1
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__A1 _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5445_ MuI._1223_ MuI._1231_ MuI._1232_ vssd1 vssd1 vccd1 vccd1 MuI._1233_ sky130_fd_sc_hd__and3_1
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1319_ AuI._0515_ vssd1 vssd1 vccd1 vccd1 AuI._0516_ sky130_fd_sc_hd__inv_2
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ _06650_ _06655_ _06649_ vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10310__B _02999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5376_ MuI._1156_ vssd1 vssd1 vccd1 vccd1 MuI._1157_ sky130_fd_sc_hd__inv_2
XFILLER_62_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07482_ _00097_ _00099_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__nor2_1
XFILLER_195_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4327_ MuI._0000_ MuI._0003_ vssd1 vssd1 vccd1 vccd1 MuI._0004_ sky130_fd_sc_hd__xnor2_1
X_09221_ _01732_ _01836_ _01835_ _01832_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__o211a_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__A1_N _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08715__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4258_ MuI._3348_ MuI._3355_ MuI._3356_ vssd1 vssd1 vccd1 vccd1 MuI._3358_ sky130_fd_sc_hd__and3_1
XANTENNA__09099__A _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _06475_ _04585_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nand2_1
XFILLER_194_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10053__A1 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ _00447_ _00449_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3556__A MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4189_ MuI._2816_ MuI._2818_ MuI._2823_ MuI._3288_ vssd1 vssd1 vccd1 vccd1 MuI._3289_
+ sky130_fd_sc_hd__o31a_1
XFILLER_148_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11250__B1 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10683__D _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _01697_ _01700_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__xor2_1
XANTENNA__10038__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0845__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _00026_ _00027_ _00146_ _00147_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__and4_1
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08731__A _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__B _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ _01860_ _01862_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__or2_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12084__A2_N _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _01231_ _01553_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nor2_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3722__C MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07509__B1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._474__A AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08867_ _01482_ _01483_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__nand3_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11019__D _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08721__A2 _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _00408_ _00409_ _00435_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a21o_1
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08798_ _02754_ _02797_ _00287_ _00267_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__and4_1
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07749_ _00365_ _00364_ _00340_ _00144_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__a211oi_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _03332_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ _01963_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10292__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10292__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _03399_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__xor2_1
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10874__C _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ _05279_ _05280_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__and3_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__B1 _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08788__A2 _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _05078_ _05082_ _05079_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11241__B1 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10595__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4907__B1 MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _04075_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__o21ai_1
XFILLER_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12292_ _04872_ _04878_ _04998_ _05133_ _04997_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__o32a_1
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5681__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5580__B1 MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ _03692_ _03693_ _03829_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__a21o_1
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1670_ AuI._0019_ AuI._0020_ AuI._0021_ vssd1 vssd1 vccd1 vccd1 AuI._0022_ sky130_fd_sc_hd__and3_1
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__B _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11544__B2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__B1 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _03927_ _03929_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__or3_1
XFILLER_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4297__A MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _03152_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__inv_2
XFILLER_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09472__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10056_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__buf_2
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3560_ MuI._1450_ MuI._1505_ vssd1 vssd1 vccd1 vccd1 MuI._1516_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11507__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13049__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07920__B1 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3491_ MuI._0339_ MuI._0746_ vssd1 vssd1 vccd1 vccd1 MuI._0757_ sky130_fd_sc_hd__and2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07423__C net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5230_ MuI.b_operand\[10\] MuI._2837_ MuI.a_operand\[6\] MuI.a_operand\[5\] vssd1
+ vssd1 vccd1 vccd1 MuI._0996_ sky130_fd_sc_hd__and4_1
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10130__B _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1104_ AuI._0240_ AuI._0243_ AuI._0223_ vssd1 vssd1 vccd1 vccd1 AuI._0314_ sky130_fd_sc_hd__mux2_1
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10958_ _03534_ _03555_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__and2_1
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5161_ MuI._0917_ MuI._0918_ MuI._0913_ vssd1 vssd1 vccd1 vccd1 MuI._0920_ sky130_fd_sc_hd__a21o_1
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1035_ AuI._0153_ AuI._0236_ AuI._0245_ AuI._0246_ vssd1 vssd1 vccd1 vccd1 AuI._0247_
+ sky130_fd_sc_hd__a31oi_1
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4112_ MuI._3197_ MuI._3210_ MuI._3211_ vssd1 vssd1 vccd1 vccd1 MuI._3212_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6060__A1 MuI._3154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _02431_ _02229_ _00783_ _05884_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nand4_1
XMuI._5092_ MuI._0795_ MuI._0843_ vssd1 vssd1 vccd1 vccd1 MuI._0844_ sky130_fd_sc_hd__or2_1
X_12628_ _00262_ _03257_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and4_1
XMuI._4043_ MuI._3066_ MuI._3069_ MuI._3140_ MuI._3141_ vssd1 vssd1 vccd1 vccd1 MuI._3143_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11599__D _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _05419_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5994_ MuI._0672_ MuI._0783_ vssd1 vssd1 vccd1 vccd1 MuI._1837_ sky130_fd_sc_hd__and2b_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4945_ MuI.a_operand\[12\] MuI.a_operand\[11\] MuI._2866_ MuI._2868_ vssd1 vssd1
+ vccd1 vccd1 MuI._0683_ sky130_fd_sc_hd__and4_1
XFILLER_99_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0819_ net118 vssd1 vssd1 vccd1 vccd1 AuI._0039_ sky130_fd_sc_hd__inv_2
XANTENNA_AuI._1252__A1 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4876_ MuI._0580_ MuI._0604_ MuI._0606_ vssd1 vssd1 vccd1 vccd1 MuI._0607_ sky130_fd_sc_hd__a21o_1
XFILLER_113_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _02096_ net116 net125 net124 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__and4_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06982_ net17 vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6615_ MuI._1290_ MuI._1457_ vssd1 vssd1 vccd1 vccd1 MuI._2520_ sky130_fd_sc_hd__nand2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3827_ MuI._2462_ MuI._2572_ vssd1 vssd1 vccd1 vccd1 MuI._2927_ sky130_fd_sc_hd__or2b_1
X_08721_ _02474_ _00030_ _00032_ _06564_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a22o_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1004__A1 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__A2 _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6546_ MuI._2426_ MuI._2443_ vssd1 vssd1 vccd1 vccd1 MuI._2444_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11417__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__C _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3758_ MuI._2847_ MuI._2848_ MuI._2857_ vssd1 vssd1 vccd1 vccd1 MuI._2858_ sky130_fd_sc_hd__nand3_1
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _01150_ _01171_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__nor2_1
XANTENNA__10321__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07603_ net119 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__buf_6
XMuI._6477_ MuI._2353_ MuI._2357_ vssd1 vssd1 vccd1 vccd1 MuI._2368_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10678__D _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3689_ MuI._2484_ vssd1 vssd1 vccd1 vccd1 MuI._2789_ sky130_fd_sc_hd__buf_2
X_08583_ _01199_ _01198_ _01192_ _01188_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__a211o_1
XFILLER_82_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5428_ MuI._1202_ MuI._1212_ MuI._1213_ vssd1 vssd1 vccd1 vccd1 MuI._1214_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4373__C MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._495__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07534_ _06488_ net129 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__nand2_1
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08467__A1 _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__B2 _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10274__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5359_ MuI._1128_ MuI._1136_ MuI._1137_ vssd1 vssd1 vccd1 vccd1 MuI._1138_ sky130_fd_sc_hd__a21bo_1
XFILLER_195_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _00082_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__buf_4
XANTENNA__10274__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__D _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _01815_ _01820_ _01816_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nand3_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07396_ _04983_ _00010_ _00013_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _01751_ _01729_ _01752_ _01434_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__o211a_1
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11774__A1 _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._469__A AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _06545_ _04649_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__nand2_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08461__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08017_ _00622_ _00633_ _00634_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__nand3_2
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10329__A2 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08611__D _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07508__C _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4117__A1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4117__B2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__inv_2
XFILLER_89_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07805__A _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _01534_ _01535_ _01536_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__nand3_2
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _02535_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__and2b_1
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10869__C _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _04742_ _04743_ _04547_ _04549_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a211oi_1
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _04515_ _04517_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nand2_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _02983_ _02980_ _04649_ _04714_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nand4_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ _04593_ _04594_ _04556_ _04466_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a211o_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10265__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _03441_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__xor2_2
XANTENNA__13261__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08355__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _02705_ _02820_ _02821_ _03306_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__a211oi_1
XFILLER_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ _03191_ _03190_ _03189_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _02865_ _05263_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
XANTENNA__11997__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13393_ _02705_ _06016_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nand2_1
XFILLER_182_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12962__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09467__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ _03497_ _05327_ _05186_ _05188_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nand4_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5553__B1 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _04975_ _05076_ _05114_ _05115_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._6300__A MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _03945_ _03946_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__nor4_1
XAuI._1653_ AuI.operand_a\[26\] AuI._0603_ vssd1 vssd1 vccd1 vccd1 AuI._0008_ sky130_fd_sc_hd__and2_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12190__A1 _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4730_ MuI._1142_ MuI._0305_ MuI._0445_ MuI._2939_ vssd1 vssd1 vccd1 vccd1 MuI._0446_
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__B2 _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07645__A1_N _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _03909_ _03910_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__o21a_1
XAuI._1584_ AuI.pe.Significand\[11\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0759_
+ sky130_fd_sc_hd__or2_1
XFILLER_96_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07137__D _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._590_ AuI.pe._131_ AuI.pe._139_ AuI.pe._144_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[11\]
+ sky130_fd_sc_hd__o21a_1
XMuI._4661_ MuI._0236_ MuI._0249_ vssd1 vssd1 vccd1 vccd1 MuI._0370_ sky130_fd_sc_hd__nor2_1
X_10108_ _02779_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__nand2_1
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11088_ _02764_ _03671_ _02350_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6400_ MuI._2107_ MuI._2244_ MuI._2282_ vssd1 vssd1 vccd1 vccd1 MuI._2283_ sky130_fd_sc_hd__and3_1
XMuI._3612_ MuI._2077_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._2088_ sky130_fd_sc_hd__nand2_1
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4592_ MuI._0292_ MuI._0293_ MuI._1263_ MuI._3246_ vssd1 vssd1 vccd1 vccd1 MuI._0294_
+ sky130_fd_sc_hd__and4bb_1
X_10039_ _02705_ _02020_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__nand2_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10141__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6331_ MuI._2205_ MuI._2206_ vssd1 vssd1 vccd1 vccd1 MuI._2207_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3543_ MuI._0339_ MuI._1318_ vssd1 vssd1 vccd1 vccd1 MuI._1329_ sky130_fd_sc_hd__and2_1
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0890__A net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3474_ MuI._0559_ vssd1 vssd1 vccd1 vccd1 MuI._0570_ sky130_fd_sc_hd__clkbuf_4
XMuI._6262_ MuI._2127_ MuI._2130_ vssd1 vssd1 vccd1 vccd1 MuI._2131_ sky130_fd_sc_hd__xnor2_2
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__A2 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__B1 _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5213_ MuI._0975_ MuI._0976_ vssd1 vssd1 vccd1 vccd1 MuI._0978_ sky130_fd_sc_hd__nand2_1
XFILLER_177_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6193_ MuI._2050_ MuI._2054_ vssd1 vssd1 vccd1 vccd1 MuI._2056_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__B _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5144_ MuI._0897_ MuI._0901_ vssd1 vssd1 vccd1 vccd1 MuI._0902_ sky130_fd_sc_hd__xnor2_1
X_07250_ _06549_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__and2b_1
XAuI._1018_ AuI._0228_ AuI._0229_ AuI._0031_ vssd1 vssd1 vccd1 vccd1 AuI._0230_ sky130_fd_sc_hd__mux2_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5075_ MuI._0795_ MuI._0825_ vssd1 vssd1 vccd1 vccd1 MuI._0826_ sky130_fd_sc_hd__and2_1
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ _06480_ _05434_ _06466_ _06479_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a22o_1
XANTENNA__12218__D _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4026_ MuI._2898_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._3126_ sky130_fd_sc_hd__nand2_1
XFILLER_185_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09096__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3553__B MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5977_ MuI._1796_ vssd1 vssd1 vccd1 vccd1 MuI._1818_ sky130_fd_sc_hd__inv_2
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4928_ MuI._0656_ MuI._0662_ MuI._0663_ vssd1 vssd1 vccd1 vccd1 MuI._0664_ sky130_fd_sc_hd__a21boi_1
X_09822_ _02424_ _02432_ _02433_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__and3_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._788_ AuI.pe._326_ AuI.pe._327_ AuI.pe._318_ vssd1 vssd1 vccd1 vccd1 AuI.pe._329_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4859_ MuI._0572_ MuI._0585_ MuI._0586_ MuI._0587_ vssd1 vssd1 vccd1 vccd1 MuI._0588_
+ sky130_fd_sc_hd__a211o_1
X_09753_ _02322_ _02395_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__nor2_1
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06965_ _05047_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08704_ _01320_ _01321_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and2_1
XFILLER_55_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09684_ _02916_ _03917_ _01918_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12372__B1_N _05218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06896_ _04305_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__buf_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6529_ MuI._2415_ MuI._2417_ MuI._2416_ MuI._2409_ vssd1 vssd1 vccd1 vccd1 MuI._2425_
+ sky130_fd_sc_hd__a211o_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08635_ _02894_ _02948_ _00267_ _00074_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__and4_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6880__A MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._468__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08566_ _01153_ _01182_ _01183_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__nor3_2
XANTENNA__08456__A _01071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10247__B2 _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _00130_ _00131_ _00134_ vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__or3_1
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08497_ _01113_ _01112_ _01048_ _01046_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__o211a_1
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07448_ _00060_ _00065_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ net39 vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__buf_4
XANTENNA__12706__A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09118_ _01711_ _01732_ _01733_ _01734_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__o211a_1
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ _02216_ _05884_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nand2_1
XANTENNA__08612__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06704__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12425__B _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3744__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09049_ _01578_ _01582_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2b_1
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09168__A2 _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12060_ _02705_ _00566_ _03306_ _02843_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a211oi_1
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12172__A1 _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _03751_ _03752_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__nand3_4
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09453__C _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ MuI.result\[21\] _02738_ _02945_ _05273_ _05852_ vssd1 vssd1 vccd1 vccd1
+ _05854_ sky130_fd_sc_hd__a221o_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input10_A a_operand[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _00281_ _02980_ _00534_ _00002_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__nand4_1
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _05778_ _05737_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nand2_1
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11844_ _04565_ _04567_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__or2_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11435__B1 _04211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11775_ _00345_ _00197_ _04575_ _04576_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__nand4_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _06545_ _03257_ _03260_ _03259_ _05959_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a32o_1
XFILLER_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07420__D _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A_N _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__inv_2
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ _03370_ _03371_ _03170_ _03172_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a211o_1
XFILLER_155_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08603__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ _06275_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__nor2_1
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ _02558_ _02560_ _02741_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08603__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5900_ MuI._1718_ MuI._1719_ MuI._1731_ MuI._1732_ vssd1 vssd1 vccd1 vccd1 MuI._1733_
+ sky130_fd_sc_hd__o211ai_1
XMuI._6880_ MuI.Exception MuI._2777_ vssd1 vssd1 vccd1 vccd1 MuI.result\[31\] sky130_fd_sc_hd__nor2_1
X_12327_ _05163_ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__and2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10136__A _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5831_ MuI._1655_ MuI._1656_ vssd1 vssd1 vccd1 vccd1 MuI._1657_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12258_ _03486_ _05262_ _05095_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__a22o_1
XFILLER_123_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._711_ AuI.pe._063_ AuI.pe._397_ AuI.pe._256_ AuI.pe._014_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._257_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._5291__D MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__A1 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5762_ MuI._1578_ MuI._1579_ MuI._1580_ vssd1 vssd1 vccd1 vccd1 MuI._1581_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._3552__A2 MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _00133_ _03099_ _05187_ _05252_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nand4_1
XFILLER_123_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1636_ AuI._0259_ AuI._0799_ AuI._0800_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[21\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12189_ _02862_ _04865_ _02722_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__o21a_1
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._642_ AuI.pe._142_ AuI.pe._053_ AuI.pe._189_ AuI.pe._192_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._193_ sky130_fd_sc_hd__a211o_1
XFILLER_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4713_ MuI._2473_ MuI._3247_ MuI._0292_ MuI._0293_ vssd1 vssd1 vccd1 vccd1 MuI._0428_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07445__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5693_ MuI._1033_ MuI._1035_ MuI._1031_ vssd1 vssd1 vccd1 vccd1 MuI._1506_ sky130_fd_sc_hd__o21bai_1
XFILLER_84_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1567_ AuI._0606_ AuI._0743_ AuI._0744_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[8\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._573_ AuI.pe._125_ AuI.pe._107_ vssd1 vssd1 vccd1 vccd1 AuI.pe._129_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4644_ MuI.a_operand\[14\] MuI._2866_ MuI._2868_ MuI.a_operand\[15\] vssd1 vssd1
+ vccd1 vccd1 MuI._0352_ sky130_fd_sc_hd__a22oi_1
XANTENNA_AuI.pe._698__A2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _02734_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[11\] sky130_fd_sc_hd__clkbuf_4
XFILLER_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1498_ AuI._0682_ AuI._0683_ vssd1 vssd1 vccd1 vccd1 AuI._0684_ sky130_fd_sc_hd__or2_2
XFILLER_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4575_ MuI._0131_ MuI._0136_ vssd1 vssd1 vccd1 vccd1 MuI._0276_ sky130_fd_sc_hd__xor2_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6254__A1 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6314_ MuI._2108_ MuI._2142_ vssd1 vssd1 vccd1 vccd1 MuI._2189_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._5844__A1_N MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3526_ MuI.b_operand\[18\] vssd1 vssd1 vccd1 vccd1 MuI._1142_ sky130_fd_sc_hd__buf_2
X_08420_ _00855_ _01036_ _01037_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__nand3_1
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09810__D net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6245_ MuI._0878_ MuI._2077_ MuI._2112_ vssd1 vssd1 vccd1 vccd1 MuI._2113_ sky130_fd_sc_hd__and3_1
XANTENNA__07180__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3829__A MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3457_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._0383_ sky130_fd_sc_hd__buf_2
XANTENNA__11426__B1 _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ _00965_ _00968_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07302_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__clkbuf_8
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6176_ MuI._1461_ MuI._1296_ MuI._1791_ MuI._1010_ vssd1 vssd1 vccd1 vccd1 MuI._2037_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3548__B MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08282_ _00866_ _00868_ _00898_ _00899_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__a211oi_4
XFILLER_177_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5127_ MuI._0865_ MuI._0881_ MuI._0882_ vssd1 vssd1 vccd1 vccd1 MuI._0883_ sky130_fd_sc_hd__nand3_2
XFILLER_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _02096_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__buf_6
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout128_A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5058_ MuI._2874_ MuI._2876_ MuI._2830_ MuI._3247_ vssd1 vssd1 vccd1 vccd1 MuI._0807_
+ sky130_fd_sc_hd__and4_1
XFILLER_192_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ _06459_ _06462_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__or3_1
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09538__C _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4009_ MuI._3107_ MuI._3108_ vssd1 vssd1 vccd1 vccd1 MuI._3109_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._3791__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _05058_ _06284_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__and2_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6297__D MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input2_A Operation[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _06544_ net115 _02454_ _02455_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4395__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07997_ _06456_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07581__A1 _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13103__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__B2 _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4826__C MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06948_ _04865_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__and3_1
X_09736_ _02380_ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__or2_1
XFILLER_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12457__A2 _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._482__A AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _02253_ _02255_ _02254_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__o21a_1
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06879_ _04122_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__buf_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13092__A _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B1 _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _01232_ _01235_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__and2b_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09598_ _02232_ _02233_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__or2b_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3739__A MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _01163_ _01161_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _02790_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__xnor2_2
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10511_ _03213_ _03214_ _03063_ _03065_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a211o_1
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _04070_ _04073_ _04071_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__o21bai_1
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5220__A2 MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13230_ _06055_ _06136_ _06101_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__or3_1
XFILLER_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _03733_ _04133_ _02969_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._5673__B MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3474__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ _05357_ _06065_ _05358_ _05749_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__or4b_1
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10373_ _00774_ _00776_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__nand2_1
XFILLER_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _04851_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__inv_2
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ _05402_ _03293_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or2b_1
XANTENNA_input58_A b_operand[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13267__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _03820_ _04736_ _04719_ _04717_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__a31o_1
XFILLER_78_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12171__A _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0948__A0 net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1421_ AuI._0140_ AuI._0252_ vssd1 vssd1 vccd1 vccd1 AuI._0607_ sky130_fd_sc_hd__or2_1
XANTENNA__07265__A _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07572__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07572__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__D _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1352_ AuI._0498_ AuI._0438_ AuI._0449_ vssd1 vssd1 vccd1 vccd1 AuI._0546_ sky130_fd_sc_hd__or3b_2
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6009__B MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10459__A1 _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11656__B1 _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B2 _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1283_ AuI._0432_ AuI._0480_ AuI._0482_ vssd1 vssd1 vccd1 vccd1 AuI._0483_ sky130_fd_sc_hd__o21ba_2
X_12945_ _05740_ _05776_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__a21o_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07324__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07324__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4360_ MuI._2055_ MuI._2852_ MuI._2873_ MuI._2875_ vssd1 vssd1 vccd1 vccd1 MuI._0040_
+ sky130_fd_sc_hd__and4_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _03110_ _05209_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nor2_1
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4291_ MuI._3325_ MuI._3337_ MuI._3332_ MuI._3336_ vssd1 vssd1 vccd1 vccd1 MuI._3391_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._3649__A MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _02752_ _04495_ _04496_ _04633_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__a31o_2
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6030_ MuI._2787_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._1876_ sky130_fd_sc_hd__nand2_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _03658_ _06613_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__nand2_1
XANTENNA__08824__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10709_ _03426_ _03427_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a21o_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__B _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ _04482_ _04483_ _04360_ _04304_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__o211a_1
XFILLER_174_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _06016_ _02825_ _06302_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__or3b_1
X_13359_ _06197_ _06252_ _06253_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__o21a_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0998_ AuI._0177_ AuI._0183_ AuI._0188_ AuI._0203_ AuI._0206_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0210_ sky130_fd_sc_hd__mux4_1
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6863_ MuI._2492_ MuI._0306_ vssd1 vssd1 vccd1 vccd1 MuI._2766_ sky130_fd_sc_hd__and2b_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5814_ MuI._1635_ MuI._1636_ MuI._1476_ vssd1 vssd1 vccd1 vccd1 MuI._1639_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3525__A2 MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _06516_ _05101_ _06517_ _06520_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22oi_1
XMuI._6794_ MuI._2643_ MuI._2696_ MuI._2698_ MuI._2700_ MuI._2716_ vssd1 vssd1 vccd1
+ vccd1 MuI._2717_ sky130_fd_sc_hd__o2111a_1
XFILLER_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12081__A _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10103__A_N _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5745_ MuI._1561_ MuI._1562_ vssd1 vssd1 vccd1 vccd1 MuI._1563_ sky130_fd_sc_hd__and2b_1
XANTENNA__07175__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1619_ AuI._0677_ AuI._0619_ AuI._0614_ vssd1 vssd1 vccd1 vccd1 AuI._0787_ sky130_fd_sc_hd__o21ai_1
X_07851_ _00465_ _00466_ _00467_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._6789__A_N MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._625_ AuI.pe._062_ AuI.pe._112_ AuI.pe._097_ AuI.pe._072_ AuI.pe._176_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._177_ sky130_fd_sc_hd__a221o_1
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06802_ _03293_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__and3_1
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5676_ MuI._1484_ MuI._1485_ MuI._1486_ vssd1 vssd1 vccd1 vccd1 MuI._1487_ sky130_fd_sc_hd__or3_1
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput2 Operation[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_4
X_07782_ _00396_ _00397_ _00399_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__nand3b_1
XANTENNA__12439__A2 _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._556_ AuI.pe._105_ AuI.pe._026_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._113_
+ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI._0898__B_N net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4627_ MuI._0187_ MuI._0186_ vssd1 vssd1 vccd1 vccd1 MuI._0333_ sky130_fd_sc_hd__nor2_1
X_09521_ _02130_ _02134_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__nand2_1
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06733_ _02550_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI.pe._540__A1 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6227__A1 MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._540__B2 AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6227__B2 MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._487_ AuI.pe._004_ vssd1 vssd1 vccd1 vccd1 AuI.pe._050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4558_ MuI._0118_ MuI._0256_ vssd1 vssd1 vccd1 vccd1 MuI._0257_ sky130_fd_sc_hd__or2_1
X_09452_ _06620_ _06437_ _02063_ _02065_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3509_ MuI._0944_ MuI._0669_ vssd1 vssd1 vccd1 vccd1 MuI._0955_ sky130_fd_sc_hd__xnor2_1
X_08403_ _06682_ _06612_ _04843_ _00000_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__a22oi_2
XANTENNA_MuI._3559__A MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4489_ MuI._0167_ MuI._0179_ MuI._0180_ vssd1 vssd1 vccd1 vccd1 MuI._0181_ sky130_fd_sc_hd__a21boi_1
X_09383_ _06593_ _04111_ _01899_ _01900_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6228_ MuI._2826_ MuI._0603_ MuI._2682_ MuI._2594_ vssd1 vssd1 vccd1 vccd1 MuI._2094_
+ sky130_fd_sc_hd__and4_1
X_08334_ _00659_ _00660_ _00588_ _00621_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a211oi_1
XANTENNA__08156__D _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08815__A1 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5196__D MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B2 _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6159_ MuI._2007_ MuI._2012_ MuI._2017_ vssd1 vssd1 vccd1 vccd1 MuI._2018_ sky130_fd_sc_hd__o21ai_1
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08265_ _02894_ _02948_ _00083_ _00098_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__and4_1
XFILLER_177_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08453__B net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07216_ _05176_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__buf_4
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ _00665_ _00813_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__and2b_1
XFILLER_119_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07147_ _03658_ _03873_ _06445_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a31o_1
XFILLER_134_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _04542_ _06067_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and2_1
XFILLER_134_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10121__B_N _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07085__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09543__A2 _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._531__A1 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _02357_ _02358_ _02362_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__nand3_1
X_10991_ _03729_ _03730_ _03548_ _03714_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__a211o_1
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07306__A1 _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__B2 _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08628__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _00231_ _00785_ _05884_ _00299_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a22o_1
XFILLER_83_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _00279_ _03424_ _00382_ _00278_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a22o_1
XFILLER_203_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11612_ _04400_ _04401_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__nor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12063__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12592_ _05453_ _05454_ _05443_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a21oi_2
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5684__A MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11543_ _04467_ _02728_ _02938_ AuI.result\[8\] vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_211_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0921_ net129 net57 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0136_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._3916__B MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._598__A1 AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ _04113_ _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__and3_1
XFILLER_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13213_ _06118_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._3755__A2 MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._098_ FuI.a_operand\[24\] FuI.a_operand\[23\] vssd1 vssd1 vccd1 vccd1 FuI._058_
+ sky130_fd_sc_hd__or2_1
XFILLER_125_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _02951_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12316__D _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0852_ AuI._0070_ net40 AuI._0071_ net9 vssd1 vssd1 vccd1 vccd1 AuI._0072_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _05953_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__inv_2
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _03045_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3860_ MuI._2418_ MuI._2958_ MuI._2959_ vssd1 vssd1 vccd1 vccd1 MuI._2960_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13075_ _05954_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__and2_1
XFILLER_2_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10287_ _03798_ _04068_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__nand2_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12026_ _04845_ _04846_ _04730_ _04734_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__o211ai_1
XMuI._3791_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._2882_ vssd1 vssd1 vccd1
+ vccd1 MuI._2891_ sky130_fd_sc_hd__o31a_1
XANTENNA_AuI._1043__B AuI._0138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5530_ MuI._1323_ MuI._1324_ MuI._1325_ vssd1 vssd1 vccd1 vccd1 MuI._1326_ sky130_fd_sc_hd__nor3b_1
XANTENNA__08742__B1 _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1404_ AuI._0579_ AuI._0588_ AuI._0591_ AuI._0587_ vssd1 vssd1 vccd1 vccd1 AuI._0593_
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._410_ AuI.pe._370_ AuI.pe._374_ AuI.pe._375_ AuI.pe._376_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._377_ sky130_fd_sc_hd__or4_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5461_ MuI._1196_ MuI._1194_ MuI._1195_ vssd1 vssd1 vccd1 vccd1 MuI._1250_ sky130_fd_sc_hd__or3_1
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1335_ AuI._0432_ AuI._0480_ AuI._0510_ AuI._0529_ vssd1 vssd1 vccd1 vccd1 AuI._0531_
+ sky130_fd_sc_hd__nor4_1
XFILLER_65_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09298__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4412_ MuI._3365_ MuI._3364_ vssd1 vssd1 vccd1 vccd1 MuI._0096_ sky130_fd_sc_hd__nor2_1
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1346__B1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5392_ MuI._0983_ MuI._0982_ MuI._0847_ vssd1 vssd1 vccd1 vccd1 MuI._1174_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07442__B _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5578__B MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1266_ net7 net122 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0467_ sky130_fd_sc_hd__mux2_2
X_12928_ _05814_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nand2_1
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4343_ MuI._0559_ MuI._3402_ MuI._0020_ MuI.a_operand\[22\] vssd1 vssd1 vccd1
+ vccd1 MuI._0022_ sky130_fd_sc_hd__a22oi_1
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1197_ AuI._0400_ AuI._0402_ vssd1 vssd1 vccd1 vccd1 AuI._0403_ sky130_fd_sc_hd__and2_1
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ _05640_ _05642_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__and2b_1
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4274_ MuI._3370_ MuI._3373_ vssd1 vssd1 vccd1 vccd1 MuI._3374_ sky130_fd_sc_hd__xnor2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6013_ MuI._1853_ MuI._1856_ vssd1 vssd1 vccd1 vccd1 MuI._1858_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12076__A _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _00483_ _00519_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__nand2_1
XFILLER_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07481__B1 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07001_ _05434_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._3746__A2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12804__A _05684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06802__A _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4938__A MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3842__A MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6846_ MuI.Exception MuI._2733_ vssd1 vssd1 vccd1 vccd1 MuI._2756_ sky130_fd_sc_hd__or2_1
XANTENNA__08720__C _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__A2 _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _03024_ _04122_ _01398_ _01397_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31o_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6777_ MuI._2683_ MuI._2697_ vssd1 vssd1 vccd1 vccd1 MuI._2698_ sky130_fd_sc_hd__xor2_1
X_07903_ _00482_ _00520_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__xnor2_2
XMuI._3989_ MuI._3060_ MuI._3061_ MuI._3063_ vssd1 vssd1 vccd1 vccd1 MuI._3089_ sky130_fd_sc_hd__and3_1
X_08883_ _01499_ _01500_ _06663_ _00033_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__and4bb_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07536__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5728_ MuI._1502_ MuI._1503_ MuI._1541_ MuI._1542_ vssd1 vssd1 vccd1 vccd1 MuI._1544_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08733__B1 _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__B1_N _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07834_ _00442_ _00450_ _00451_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__nand3_1
XFILLER_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI.pe._608_ AuI.pe._125_ AuI.pe._050_ AuI.pe._078_ AuI.pe._089_ AuI.pe._160_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._161_ sky130_fd_sc_hd__a221o_1
XANTENNA__10978__B _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5659_ MuI._1318_ MuI._1813_ MuI._0246_ MuI._0420_ vssd1 vssd1 vccd1 vccd1 MuI._1468_
+ sky130_fd_sc_hd__nand4_1
XFILLER_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07765_ _06544_ _00382_ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__nand2_1
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._539_ AuI.pe._096_ vssd1 vssd1 vccd1 vccd1 AuI.pe._097_ sky130_fd_sc_hd__buf_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11155__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09504_ _01891_ _01988_ _01987_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__o21ai_1
X_06716_ net108 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__clkbuf_8
XFILLER_65_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07839__A2 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ _00305_ _00307_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ _06663_ _06433_ _02055_ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__and4_1
XANTENNA__10843__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10843__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13370__A _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _01983_ _01892_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5000__C MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08317_ _00909_ _00932_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _01808_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__xor2_1
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _00863_ _00864_ _00865_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__a21o_2
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0863__A2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08196__A_N _00665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _00795_ _00796_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__xor2_2
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10210_ _02891_ _02860_ _02859_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _03781_ _03784_ _03782_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o21bai_1
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09726__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06712__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08630__C _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _03755_ _05906_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._6151__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._752__A1 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_AuI.pe._752__B2 AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A2_N _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12520__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10888__B _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__A _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1120_ AuI._0328_ AuI._0326_ vssd1 vssd1 vccd1 vccd1 AuI._0329_ sky130_fd_sc_hd__nor2_2
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _03363_ _03367_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a211oi_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08077__C _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ _02744_ _03974_ _02944_ _05058_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a22o_1
XAuI._1051_ AuI._0150_ AuI._0151_ vssd1 vssd1 vccd1 vccd1 AuI._0262_ sky130_fd_sc_hd__and2_2
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ _05440_ _05322_ _05458_ _05459_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a211oi_1
XFILLER_169_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _00502_ _05123_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10062__A2 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _04307_ _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__or2_1
XFILLER_184_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0904_ AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0124_ sky130_fd_sc_hd__clkbuf_4
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _02840_ _05649_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nand2_1
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0877__B net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__B _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4961_ MuI._0697_ MuI._0699_ vssd1 vssd1 vccd1 vccd1 MuI._0700_ sky130_fd_sc_hd__and2b_1
X_10408_ _00749_ _00803_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__a21oi_1
XAuI._0835_ AuI._0053_ net34 AuI._0054_ net123 vssd1 vssd1 vccd1 vccd1 AuI._0055_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output89_A net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11388_ _02935_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4758__A MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6700_ MuI._2603_ MuI._2383_ vssd1 vssd1 vccd1 vccd1 MuI._2613_ sky130_fd_sc_hd__and2b_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3912_ MuI._2817_ MuI._2787_ MuI._2941_ vssd1 vssd1 vccd1 vccd1 MuI._3012_ sky130_fd_sc_hd__and3_1
XFILLER_113_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08540__C _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4892_ MuI._0622_ MuI._0623_ MuI._1263_ MuI._0445_ vssd1 vssd1 vccd1 vccd1 MuI._0624_
+ sky130_fd_sc_hd__and4bb_1
X_10339_ _00734_ _00736_ _00735_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__o21bai_1
XFILLER_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13127_ _05961_ _05964_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a21o_1
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6631_ MuI._1460_ MuI._1645_ MuI._1764_ vssd1 vssd1 vccd1 vccd1 MuI._2537_ sky130_fd_sc_hd__o21a_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3843_ MuI._2941_ MuI._2942_ vssd1 vssd1 vccd1 vccd1 MuI._2943_ sky130_fd_sc_hd__xnor2_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _03669_ _05585_ _05887_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4908__D MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0893__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6562_ MuI._2452_ MuI._2454_ vssd1 vssd1 vccd1 vccd1 MuI._2461_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ net61 _04800_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nand2_1
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3774_ MuI._2873_ vssd1 vssd1 vccd1 vccd1 MuI._2874_ sky130_fd_sc_hd__clkbuf_4
XFILLER_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1031__A2 net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5513_ MuI._0100_ MuI._3262_ MuI.a_operand\[4\] MuI._0020_ vssd1 vssd1 vccd1
+ vccd1 MuI._1308_ sky130_fd_sc_hd__and4_1
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6493_ MuI._0793_ MuI._1841_ MuI._2005_ MuI._2367_ MuI._2384_ vssd1 vssd1 vccd1
+ vccd1 MuI._2386_ sky130_fd_sc_hd__a2111o_1
XFILLER_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13067__A2 _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5444_ MuI._1166_ MuI._1228_ MuI._1217_ MuI._1227_ vssd1 vssd1 vccd1 vccd1 MuI._1232_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07550_ _00158_ _00159_ _00167_ vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__nand3_1
XAuI._1318_ AuI._0438_ AuI._0408_ AuI._0421_ AuI._0514_ vssd1 vssd1 vccd1 vccd1 AuI._0515_
+ sky130_fd_sc_hd__o211a_2
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5375_ MuI._1139_ MuI._1152_ MuI._1154_ MuI._1155_ vssd1 vssd1 vccd1 vccd1 MuI._1156_
+ sky130_fd_sc_hd__a211o_1
X_07481_ _03099_ _00098_ _00047_ _03056_ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__a22oi_1
XAuI._1249_ AuI._0389_ AuI._0449_ AuI._0450_ vssd1 vssd1 vccd1 vccd1 AuI._0451_ sky130_fd_sc_hd__o21ai_4
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4326_ MuI._0001_ MuI._0002_ vssd1 vssd1 vccd1 vccd1 MuI._0003_ sky130_fd_sc_hd__nor2_1
X_09220_ _01798_ _01799_ _01807_ _01808_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__o22a_1
XFILLER_195_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4613__B1 MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4257_ MuI._3348_ MuI._3355_ MuI._3356_ vssd1 vssd1 vccd1 vccd1 MuI._3357_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08715__C _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ _00162_ _04638_ _00033_ _00164_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22oi_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10319__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _00717_ _00718_ _00714_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__a21o_1
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4188_ MuI._2824_ MuI._2832_ vssd1 vssd1 vccd1 vccd1 MuI._3288_ sky130_fd_sc_hd__nand2_1
XANTENNA__10053__A2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _01698_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11250__B2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10038__B _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _00026_ _00027_ _00146_ _00147_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__a22oi_2
XFILLER_190_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout110_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 b_operand[30] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_4
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08731__B _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10980__C _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6118__B1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09984_ _02646_ _01865_ _02648_ _02649_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a211oi_4
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6829_ MuI._2746_ vssd1 vssd1 vccd1 vccd1 MuI.result\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09843__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _06620_ _00036_ _01229_ _01230_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07509__A1 _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07509__B2 _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13365__A _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08866_ _01283_ _01282_ _01281_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__o21ai_1
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07363__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07817_ _00433_ _00434_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__and2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _01365_ _01381_ _01413_ _01414_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a211oi_4
XANTENNA__09281__C _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._498__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07748_ _00144_ _00340_ _00364_ _00365_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__o211a_1
XANTENNA_MuI._3655__B2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _00285_ _00296_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__xnor2_2
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11613__A _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09418_ _01964_ _02037_ _01959_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10292__A2 _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__and2b_1
XFILLER_40_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07693__B1 _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__A _00810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10874__D _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _06479_ _06480_ _00084_ _04574_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and4_1
XANTENNA__09434__A1 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10229__A _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__B2 _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _05205_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4907__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ _04075_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._4907__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _04999_ _04996_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nor2_1
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11242_ _04001_ _04003_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._5681__B MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13259__B _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11544__A2 _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12741__B2 _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _06680_ _00163_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3913__C MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10124_ _02798_ _02799_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nor2_2
XANTENNA_input40_A b_operand[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0917__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10055_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09472__B _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13049__A2 _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__C _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._489__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07920__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3490_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._0746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07423__D _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1103_ AuI._0177_ AuI._0310_ AuI._0311_ AuI._0312_ AuI._0233_ AuI._0307_ vssd1
+ vssd1 vccd1 vccd1 AuI._0313_ sky130_fd_sc_hd__mux4_1
X_10957_ _03514_ _03557_ _03695_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__a21o_2
XFILLER_73_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5160_ MuI._0913_ MuI._0917_ MuI._0918_ vssd1 vssd1 vccd1 vccd1 MuI._0919_ sky130_fd_sc_hd__nand3_1
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1034_ AuI._0157_ AuI._0211_ vssd1 vssd1 vccd1 vccd1 AuI._0246_ sky130_fd_sc_hd__and2_1
XANTENNA__07684__B1 _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11480__B2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4111_ MuI._2864_ MuI._3196_ MuI._3182_ vssd1 vssd1 vccd1 vccd1 MuI._3211_ sky130_fd_sc_hd__nand3_1
X_10888_ _02528_ _03247_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nand2_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3657__A MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5091_ MuI._0828_ MuI._0842_ vssd1 vssd1 vccd1 vccd1 MuI._0843_ sky130_fd_sc_hd__nor2_1
XFILLER_176_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12627_ _00921_ _01206_ _03444_ _05948_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__and4_1
XANTENNA__10139__A _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4042_ MuI._3066_ MuI._3069_ MuI._3140_ MuI._3141_ vssd1 vssd1 vccd1 vccd1 MuI._3142_
+ sky130_fd_sc_hd__nand4_1
XFILLER_157_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12558_ _05399_ _05287_ _05418_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand3_1
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12980__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11509_ _04088_ _04090_ _04289_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__o211ai_4
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ _05266_ _05236_ _05344_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__o211a_1
XFILLER_172_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5993_ MuI._1766_ MuI._1816_ MuI._1830_ MuI._1834_ vssd1 vssd1 vccd1 vccd1 MuI._1836_
+ sky130_fd_sc_hd__o31a_2
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4944_ MuI._0674_ MuI._0678_ MuI._0681_ vssd1 vssd1 vccd1 vccd1 MuI._0682_ sky130_fd_sc_hd__o21ai_1
XFILLER_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0818_ net117 vssd1 vssd1 vccd1 vccd1 AuI._0038_ sky130_fd_sc_hd__inv_2
XFILLER_140_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4875_ MuI._0489_ MuI._0605_ vssd1 vssd1 vccd1 vccd1 MuI._0606_ sky130_fd_sc_hd__or2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _05220_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[19\] sky130_fd_sc_hd__buf_2
XFILLER_140_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6614_ MuI._1290_ MuI._1457_ vssd1 vssd1 vccd1 vccd1 MuI._2519_ sky130_fd_sc_hd__or2_1
XFILLER_140_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3826_ MuI._2865_ MuI._2924_ MuI._2925_ vssd1 vssd1 vccd1 vccd1 MuI._2926_ sky130_fd_sc_hd__a21oi_2
XANTENNA_AuI._1512__A AuI._0116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _06564_ _02474_ _00030_ _00032_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3885__A1 MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3885__B2 MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__A _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6545_ MuI._2438_ MuI._2442_ vssd1 vssd1 vccd1 vccd1 MuI._2443_ sky130_fd_sc_hd__nand2_1
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3757_ MuI._2849_ MuI._2851_ MuI._2855_ MuI._2856_ vssd1 vssd1 vccd1 vccd1 MuI._2857_
+ sky130_fd_sc_hd__a31o_1
X_08651_ _01263_ _01267_ _01245_ _01268_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__a211oi_2
XFILLER_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11417__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10321__B _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07602_ _03013_ _06613_ _00218_ _00219_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__nand4_1
XFILLER_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6476_ MuI._2307_ MuI._2339_ MuI._2366_ vssd1 vssd1 vccd1 vccd1 MuI._2367_ sky130_fd_sc_hd__or3_1
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3688_ MuI._2550_ MuI._2517_ MuI._2495_ MuI._2773_ vssd1 vssd1 vccd1 vccd1 MuI._2788_
+ sky130_fd_sc_hd__and4_1
X_08582_ _01188_ _01192_ _01198_ _01199_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__o211ai_4
XFILLER_208_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5427_ MuI._1184_ MuI._1185_ MuI._1201_ vssd1 vssd1 vccd1 vccd1 MuI._1213_ sky130_fd_sc_hd__a21o_1
XANTENNA__07911__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ _06494_ _00150_ net128 net28 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._4373__D MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__B2 _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__A2 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08726__B _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5358_ MuI._1129_ MuI._1130_ MuI._1135_ vssd1 vssd1 vccd1 vccd1 MuI._1137_ sky130_fd_sc_hd__nand3_1
XFILLER_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11433__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07464_ net35 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__buf_2
XANTENNA__10274__A2 _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4309_ MuI._3263_ MuI._3269_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._3409_ sky130_fd_sc_hd__and3b_1
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _01815_ _01816_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21o_1
XMuI._5289_ MuI._0984_ MuI._1060_ vssd1 vssd1 vccd1 vccd1 MuI._1061_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07395_ _00011_ _06591_ _05036_ _00012_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__a22o_1
XFILLER_176_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13346__B1_N _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ _01431_ _01432_ _01433_ _01408_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11774__A2 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ _01681_ _01682_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__and2b_1
XFILLER_190_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08461__B _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08016_ _06508_ _06498_ _06507_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__a21o_1
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4117__A2 MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _01676_ _01767_ _01844_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__nand3b_2
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08918_ _01288_ _01285_ _01287_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a21o_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _02259_ _03917_ _02534_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a21o_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07093__A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__D _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _01455_ _01460_ _01456_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__nand3_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _04666_ _04667_ _04663_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a21o_1
XFILLER_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _03443_ _04649_ _00040_ _00281_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a22o_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _04556_ _04466_ _04593_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__o211ai_4
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09655__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10265__A2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ _03463_ _03464_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__nand2_1
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13461_ _01330_ _06374_ _06375_ _02741_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__o211a_2
X_10673_ _03388_ _03386_ _03387_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__nand3_1
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12412_ _05261_ _02899_ _04635_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__mux2_1
XANTENNA__09958__A2 _02584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13392_ _01322_ _06304_ _02699_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__or3_4
XANTENNA__08652__A _01150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6220__A1_N MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12962__B2 _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__B _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _03497_ _05327_ _05186_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a22o_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__B _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5553__A1 MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12274_ _05111_ _05113_ _05077_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o21a_1
XFILLER_181_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6300__B MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12714__B2 _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _03983_ _03984_ _03754_ _03947_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__o211a_1
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1652_ AuI.exponent_sub\[3\] AuI._0769_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0007_
+ sky130_fd_sc_hd__o21a_1
XFILLER_107_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12902__A _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__A2 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _02539_ _05895_ _05959_ _02496_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__a22o_1
XAuI._1583_ AuI._0693_ AuI._0750_ AuI._0757_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0758_
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06900__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3940__A MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4660_ MuI._0326_ MuI._0367_ MuI._0368_ vssd1 vssd1 vccd1 vccd1 MuI._0369_ sky130_fd_sc_hd__a21o_1
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _02780_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__nor2b_2
XFILLER_49_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11087_ _02565_ _03836_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__nor2_1
XANTENNA__08099__A _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3611_ MuI._2066_ vssd1 vssd1 vccd1 vccd1 MuI._2077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4591_ MuI._1802_ MuI._2319_ MuI._0101_ MuI._1307_ vssd1 vssd1 vccd1 vccd1 MuI._0293_
+ sky130_fd_sc_hd__a22oi_1
X_10038_ _02705_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__nand2_1
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10141__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6028__A MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6330_ MuI._2077_ MuI._2120_ MuI._2180_ MuI._2181_ vssd1 vssd1 vccd1 vccd1 MuI._2206_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3542_ MuI._1307_ vssd1 vssd1 vccd1 vccd1 MuI._1318_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._0890__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6261_ MuI._2128_ MuI._2129_ vssd1 vssd1 vccd1 vccd1 MuI._2130_ sky130_fd_sc_hd__nor2_1
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3473_ MuI.a_operand\[21\] vssd1 vssd1 vccd1 vccd1 MuI._0559_ sky130_fd_sc_hd__clkbuf_4
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__A1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5212_ MuI._0973_ MuI._0974_ MuI._0969_ MuI._0972_ vssd1 vssd1 vccd1 vccd1 MuI._0976_
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__09646__B2 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _04675_ _04695_ _04806_ _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__a211o_1
XFILLER_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6192_ MuI._2051_ MuI._2053_ vssd1 vssd1 vccd1 vccd1 MuI._2054_ sky130_fd_sc_hd__nor2_1
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5586__B MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5143_ MuI._0898_ MuI._0899_ vssd1 vssd1 vccd1 vccd1 MuI._0901_ sky130_fd_sc_hd__nor2_1
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08265__C _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1017_ net68 net36 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0229_ sky130_fd_sc_hd__mux2_1
XFILLER_177_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5074_ MuI._2919_ MuI._0315_ MuI.a_operand\[0\] MuI._2800_ vssd1 vssd1 vccd1
+ vccd1 MuI._0825_ sky130_fd_sc_hd__a22o_1
XANTENNA__09658__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _06479_ _06480_ net20 _06466_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__and4_1
XFILLER_185_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4025_ MuI._3123_ MuI._3124_ vssd1 vssd1 vccd1 vccd1 MuI._3125_ sky130_fd_sc_hd__nor2_1
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11756__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5544__A1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07178__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09096__C net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5976_ MuI._0740_ MuI._0778_ vssd1 vssd1 vccd1 vccd1 MuI._1817_ sky130_fd_sc_hd__xnor2_4
XANTENNA_MuI._3553__C MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4927_ MuI._0654_ MuI._0655_ vssd1 vssd1 vccd1 vccd1 MuI._0663_ sky130_fd_sc_hd__nand2_1
XANTENNA__12181__A2 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _02467_ _02471_ _02472_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__or3_1
XFILLER_113_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06810__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._787_ AuI.pe._318_ AuI.pe._326_ AuI.pe._327_ vssd1 vssd1 vccd1 vccd1 AuI.pe._328_
+ sky130_fd_sc_hd__and3_1
XFILLER_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4858_ MuI._0517_ MuI._0518_ MuI._0519_ vssd1 vssd1 vccd1 vccd1 MuI._0587_ sky130_fd_sc_hd__and3_1
XFILLER_140_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ _02324_ _02346_ _02398_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__o21bai_1
X_06964_ _05036_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__buf_4
XANTENNA__10332__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3809_ MuI._1472_ MuI._2844_ MuI._2845_ MuI._1010_ vssd1 vssd1 vccd1 vccd1 MuI._2909_
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08703_ _01200_ _01201_ _01319_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__a21o_1
XMuI._4789_ MuI._0507_ MuI._0509_ vssd1 vssd1 vccd1 vccd1 MuI._0511_ sky130_fd_sc_hd__xnor2_1
X_09683_ _02090_ _02163_ _02161_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a21boi_1
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06895_ _04294_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__buf_4
XFILLER_55_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6528_ MuI._2421_ MuI._2423_ vssd1 vssd1 vccd1 vccd1 MuI._2424_ sky130_fd_sc_hd__nand2_1
XFILLER_67_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _01249_ _01251_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__or2b_1
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6459_ MuI._2346_ MuI._2347_ vssd1 vssd1 vccd1 vccd1 MuI._2348_ sky130_fd_sc_hd__or2b_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07641__A _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _01129_ _01131_ _01181_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__nor3_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12259__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10247__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07516_ _00132_ _00047_ _00048_ _00133_ vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__a22oi_2
X_08496_ _01046_ _01048_ _01112_ _01113_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__a211oi_2
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ _00061_ _00064_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__nor2_1
XFILLER_196_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07378_ _06628_ _06635_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and2_1
XFILLER_164_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12706__B _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09117_ _01711_ _01732_ _01733_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__o211ai_2
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__A2 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12425__C _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ _01664_ _01663_ _01590_ _01566_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__a211oi_1
XFILLER_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _03567_ _03566_ _03565_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__a21bo_1
XFILLER_78_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06720__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3760__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10242__A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A1 _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__D _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12961_ _05338_ _02727_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A1 _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _03443_ _05112_ _06525_ _00290_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a22o_1
XFILLER_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _05653_ _05734_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__or2b_1
XFILLER_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04644_ _04646_ _04650_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or3_1
XFILLER_45_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12176__A1_N _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _00283_ _00197_ _04575_ _04576_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__a22o_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08085__C _00702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _03248_ _03251_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__nand2_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._616__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13188__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11801__A _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13444_ _06296_ _06328_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__or2_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _03170_ _03172_ _03370_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o211ai_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1327__A AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10587_ _03294_ _03297_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__or2_1
XANTENNA__08603__A2 _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ _06286_ _06287_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__nand2_1
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12326_ _05168_ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__xor2_1
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10136__B _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5830_ MuI._0718_ MuI._0717_ vssd1 vssd1 vccd1 vccd1 MuI._1656_ sky130_fd_sc_hd__and2b_1
XFILLER_182_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6030__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _02983_ _02984_ _03047_ _06477_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nand4_1
XANTENNA__12699__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._710_ AuI.pe.significand\[3\] AuI.pe._394_ AuI.pe._395_ AuI.pe._255_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._256_ sky130_fd_sc_hd__and4_1
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5761_ MuI._1484_ MuI._1486_ MuI._1485_ vssd1 vssd1 vccd1 vccd1 MuI._1580_ sky130_fd_sc_hd__o21bai_1
XANTENNA_output71_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1635_ AuI.pe.Significand\[21\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0800_
+ sky130_fd_sc_hd__or2_1
X_11208_ _00081_ _05187_ _05252_ _00086_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a22o_1
X_12188_ _02402_ _05008_ _05007_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__and3_1
XFILLER_122_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._641_ AuI.pe._071_ AuI.pe._391_ AuI.pe._041_ AuI.pe._158_ AuI.pe._191_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._192_ sky130_fd_sc_hd__a221o_1
XMuI._4712_ MuI._0423_ MuI._0425_ vssd1 vssd1 vccd1 vccd1 MuI._0426_ sky130_fd_sc_hd__nor2_1
XFILLER_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5692_ MuI._1029_ MuI._1048_ MuI._1049_ vssd1 vssd1 vccd1 vccd1 MuI._1504_ sky130_fd_sc_hd__nand3_1
XANTENNA__11248__A _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1566_ AuI.pe.Significand\[8\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0744_
+ sky130_fd_sc_hd__or2_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _03890_ _03888_ _03889_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nand3_2
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._572_ AuI.pe._084_ AuI.pe._050_ AuI.pe._079_ AuI.pe._059_ AuI.pe._127_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._128_ sky130_fd_sc_hd__a221o_1
XMuI._4643_ MuI._2440_ MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 MuI._0351_ sky130_fd_sc_hd__nand2_1
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1497_ AuI._0564_ AuI._0566_ vssd1 vssd1 vccd1 vccd1 AuI._0683_ sky130_fd_sc_hd__nor2_1
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4574_ MuI._0266_ MuI._0272_ MuI._0274_ vssd1 vssd1 vccd1 vccd1 MuI._0275_ sky130_fd_sc_hd__a21o_1
XFILLER_92_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6313_ MuI._2185_ MuI._2186_ vssd1 vssd1 vccd1 vccd1 MuI._2188_ sky130_fd_sc_hd__nand2_1
XMuI._3525_ MuI._0889_ MuI._0537_ MuI._0757_ MuI._1120_ vssd1 vssd1 vccd1 vccd1 MuI._1131_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6244_ MuI._2109_ MuI._2111_ vssd1 vssd1 vccd1 vccd1 MuI._2112_ sky130_fd_sc_hd__nor2_1
XFILLER_211_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3456_ MuI._0361_ vssd1 vssd1 vccd1 vccd1 MuI._0372_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07180__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _00966_ _00967_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__nor2_1
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11426__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3829__B MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07301_ net10 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__buf_4
XMuI._6175_ MuI.b_operand\[17\] MuI._2843_ vssd1 vssd1 vccd1 vccd1 MuI._2036_ sky130_fd_sc_hd__nand2_1
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ _00580_ _00581_ _00583_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__nor3_2
XANTENNA__12807__A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5126_ MuI._0879_ MuI._0880_ MuI._0871_ vssd1 vssd1 vccd1 vccd1 MuI._0882_ sky130_fd_sc_hd__a21o_1
XANTENNA__13402__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ _06511_ _06512_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__nand3_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06805__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5057_ MuI._0799_ MuI._0805_ vssd1 vssd1 vccd1 vccd1 MuI._0806_ sky130_fd_sc_hd__or2b_1
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07163_ _06463_ _05627_ net130 _02107_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a22oi_2
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4008_ MuI._2817_ MuI._2789_ vssd1 vssd1 vccd1 vccd1 MuI._3108_ sky130_fd_sc_hd__nand2_1
XANTENNA__09538__D _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10182__A_N _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3791__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ _06410_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6190__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6190__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13351__A1 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5959_ MuI._1796_ MuI._1797_ vssd1 vssd1 vccd1 vccd1 MuI._1798_ sky130_fd_sc_hd__and2_1
XANTENNA__13351__B2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _02454_ _02455_ _06544_ net115 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__and4bb_1
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11158__A _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07996_ _00602_ _00612_ _00613_ _00317_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__o211ai_4
XANTENNA_MuI._4395__B MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13103__B2 _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__A2 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4826__D MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _02604_ _03917_ _02378_ _02379_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a211oi_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06947_ _04854_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07869__B1 _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _02304_ _02305_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__nand3_2
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06878_ _04111_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__buf_4
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08530__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _01233_ _01234_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__xnor2_2
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09597_ _02222_ _02225_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__xor2_1
XANTENNA__13406__A2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3739__B MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _01149_ _01165_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__nor2_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08294__B1 _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ _00923_ _00922_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__nor2_1
XFILLER_211_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ _03063_ _03065_ _03213_ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__o211ai_1
XFILLER_211_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11490_ _04074_ _04083_ _04082_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__a21o_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10441_ _02968_ _02967_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__or2b_1
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10372_ _03065_ _03066_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__nor2_1
X_13160_ _05919_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__or2_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12111_ _04810_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__xor2_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13091_ _05988_ _05989_ _03134_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__o21a_1
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__B1 _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _04862_ _04863_ _04751_ _04753_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a211o_2
XANTENNA__07546__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13267__B _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4586__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3490__A MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1420_ AuI._0258_ vssd1 vssd1 vccd1 vccd1 AuI._0606_ sky130_fd_sc_hd__buf_2
XANTENNA_AuI._0948__A1 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07265__B _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07572__A2 _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1351_ AuI._0536_ AuI._0545_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[17\]
+ sky130_fd_sc_hd__xor2_2
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09761__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11656__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__A2 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12944_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nand2_1
XAuI._1282_ AuI._0458_ AuI._0479_ AuI._0481_ AuI._0469_ vssd1 vssd1 vccd1 vccd1 AuI._0482_
+ sky130_fd_sc_hd__a22o_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__A2 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07281__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08808__C _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _03974_ _03973_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__nor2_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4290_ MuI._3389_ MuI._3379_ vssd1 vssd1 vccd1 vccd1 MuI._3390_ sky130_fd_sc_hd__xnor2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _04619_ _04621_ _04623_ _03315_ _04632_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__a221o_1
XFILLER_61_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11757_ _00550_ _04557_ _04558_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21bo_2
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12627__A _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08824__B net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ _06680_ _00398_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__inv_2
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3665__A MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _02815_ _06302_ _06334_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__a21o_1
XANTENNA__13030__B1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10639_ _03798_ _04197_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__nand2_1
XFILLER_155_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _06196_ _06252_ _06253_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__o21a_1
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0896__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0997_ AuI._0208_ vssd1 vssd1 vccd1 vccd1 AuI._0209_ sky130_fd_sc_hd__buf_2
XFILLER_170_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6862_ MuI._2735_ MuI._2764_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[24\]
+ sky130_fd_sc_hd__a21oi_1
X_12309_ _03013_ _05895_ _05959_ _02970_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a22o_1
X_13289_ _06196_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__nand2_1
XFILLER_170_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5813_ MuI._1476_ MuI._1635_ MuI._1636_ vssd1 vssd1 vccd1 vccd1 MuI._1638_ sky130_fd_sc_hd__and3_1
XFILLER_170_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6793_ MuI._2683_ MuI._2701_ MuI._2702_ MuI._2705_ MuI._2714_ vssd1 vssd1 vccd1
+ vccd1 MuI._2716_ sky130_fd_sc_hd__o2111a_1
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07456__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12081__B _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5744_ MuI._2754_ MuI._0110_ MuI.a_operand\[1\] MuI._1307_ vssd1 vssd1 vccd1
+ vccd1 MuI._1562_ sky130_fd_sc_hd__a22o_1
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1618_ AuI._0259_ AuI._0785_ AuI._0786_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[17\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07850_ _00465_ _00466_ _00467_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__and3_1
XAuI.pe._624_ AuI.pe.significand\[4\] AuI.pe._119_ vssd1 vssd1 vccd1 vccd1 AuI.pe._176_
+ sky130_fd_sc_hd__and2_1
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5675_ MuI._2845_ MuI._0088_ MuI._2319_ MuI._2844_ vssd1 vssd1 vccd1 vccd1 MuI._1486_
+ sky130_fd_sc_hd__a22oi_2
X_06801_ _03282_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__buf_4
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1549_ AuI.pe.Significand\[5\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0730_
+ sky130_fd_sc_hd__or2_1
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07781_ _06565_ _02485_ _00398_ _05563_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__nand4_1
XFILLER_83_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput3 Operation[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09103__A1_N _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4626_ MuI._0329_ MuI._0331_ vssd1 vssd1 vccd1 vccd1 MuI._0332_ sky130_fd_sc_hd__nor2_1
XAuI.pe._555_ AuI.pe._391_ vssd1 vssd1 vccd1 vccd1 AuI.pe._112_ sky130_fd_sc_hd__buf_2
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09520_ _02131_ _02133_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__or2b_1
X_06732_ _02539_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__buf_8
XFILLER_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI.pe._540__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6227__A2 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._486_ AuI.pe._048_ vssd1 vssd1 vccd1 vccd1 AuI.pe._049_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07191__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4557_ MuI._0094_ MuI._0095_ MuI._0117_ vssd1 vssd1 vccd1 vccd1 MuI._0256_ sky130_fd_sc_hd__o21a_1
XFILLER_80_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ _02052_ _02060_ _02073_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a21oi_2
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3508_ MuI._0592_ MuI._0471_ vssd1 vssd1 vccd1 vccd1 MuI._0944_ sky130_fd_sc_hd__nand2_1
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08402_ _06593_ _04714_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__nand2_1
XMuI._4488_ MuI._0164_ MuI._0166_ vssd1 vssd1 vccd1 vccd1 MuI._0180_ sky130_fd_sc_hd__or2b_1
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3559__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ _01997_ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__nor2_1
XFILLER_178_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6227_ MuI._0603_ MuI._2914_ MuI._2594_ MuI._2826_ vssd1 vssd1 vccd1 vccd1 MuI._2093_
+ sky130_fd_sc_hd__a22oi_1
XMuI._3439_ MuI.a_operand\[28\] MuI.b_operand\[28\] vssd1 vssd1 vccd1 vccd1 MuI._0185_
+ sky130_fd_sc_hd__or2_1
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _00947_ _00950_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__or2_2
XANTENNA__08595__A_N _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A2 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6158_ MuI._2013_ MuI._2016_ vssd1 vssd1 vccd1 vccd1 MuI._2017_ sky130_fd_sc_hd__xnor2_1
X_08264_ _00574_ _00880_ _00881_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__nand3_1
XFILLER_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5109_ MuI._0859_ MuI._0862_ vssd1 vssd1 vccd1 vccd1 MuI._0863_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08453__C _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6089_ MuI._1939_ MuI._1940_ vssd1 vssd1 vccd1 vccd1 MuI._1941_ sky130_fd_sc_hd__nand2_1
X_07215_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__buf_4
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ _00666_ _00812_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__xor2_1
XFILLER_192_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10057__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09776__B1 _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _06444_ _06442_ _03960_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__and4_1
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07077_ _06243_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13324__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07366__A _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4974__A2_N MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ _00593_ _00596_ vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__and2b_1
XFILLER_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1430__A AuI._0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _02357_ _02358_ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a21o_1
XANTENNA__11616__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._531__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _03548_ _03714_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__o211ai_2
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07306__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08628__C _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _02258_ _02262_ _02261_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a21o_1
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _05400_ _05404_ _05401_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__o21bai_1
XFILLER_70_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11611_ _00124_ _00125_ _06525_ _05252_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__and4_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08267__B1 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _05443_ _05453_ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__and3_2
XFILLER_169_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10074__B1 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5684__B MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3485__A MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0920_ AuI._0135_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[27\] sky130_fd_sc_hd__buf_2
X_11473_ _04131_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__inv_2
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._097_ FuI._052_ FuI._057_ FuI.a_operand\[8\] vssd1 vssd1 vccd1 vccd1 FuI._020_
+ sky130_fd_sc_hd__o21a_1
X_13212_ _06026_ _06027_ _06024_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ _03122_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__and2b_1
XAuI._0851_ net41 vssd1 vssd1 vccd1 vccd1 AuI._0071_ sky130_fd_sc_hd__inv_2
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13143_ _06035_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__xor2_1
XFILLER_125_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10355_ _03046_ _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _05971_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2_1
X_10286_ _02973_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nor2_2
XFILLER_140_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3790_ MuI.a_operand\[24\] MuI.a_operand\[23\] MuI.a_operand\[26\] vssd1 vssd1
+ vccd1 vccd1 MuI._2890_ sky130_fd_sc_hd__or3_4
X_12025_ _04730_ _04734_ _04845_ _04846_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__a211o_1
XFILLER_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1403_ AuI._0589_ AuI._0592_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[22\]
+ sky130_fd_sc_hd__xor2_4
XANTENNA__10133__C _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__A1 _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08742__B2 _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5460_ MuI._1247_ MuI._1248_ vssd1 vssd1 vccd1 vccd1 MuI._1249_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1334_ AuI._0510_ AuI._0529_ vssd1 vssd1 vccd1 vccd1 AuI._0530_ sky130_fd_sc_hd__nor2_1
XFILLER_207_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4411_ MuI._0084_ MuI._0092_ MuI._0093_ vssd1 vssd1 vccd1 vccd1 MuI._0095_ sky130_fd_sc_hd__and3_1
XANTENNA__09641__D _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__A2 _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5391_ MuI._0983_ MuI._0847_ MuI._0982_ vssd1 vssd1 vccd1 vccd1 MuI._1173_ sky130_fd_sc_hd__and3_1
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1265_ AuI._0420_ AuI._0465_ vssd1 vssd1 vccd1 vccd1 AuI._0466_ sky130_fd_sc_hd__nand2_1
X_12927_ _03744_ _05391_ _05722_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nand3_1
XFILLER_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4342_ MuI._0018_ vssd1 vssd1 vccd1 vccd1 MuI._0020_ sky130_fd_sc_hd__clkbuf_4
XFILLER_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1196_ AuI._0362_ AuI._0401_ AuI._0380_ vssd1 vssd1 vccd1 vccd1 AuI._0402_ sky130_fd_sc_hd__o21ai_1
X_12858_ _05740_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__and2_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4273_ MuI._3372_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._3373_ sky130_fd_sc_hd__nand2_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08258__B1 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ _04312_ _04487_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nand2_1
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6012_ MuI._1854_ MuI._1855_ vssd1 vssd1 vccd1 vccd1 MuI._1856_ sky130_fd_sc_hd__nor2_1
XANTENNA__12357__A _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12789_ _05565_ _05570_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08554__B _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07481__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07481__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07000_ net20 vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__clkbuf_4
XFILLER_179_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11565__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4938__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13306__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6845_ MuI._2755_ vssd1 vssd1 vccd1 vccd1 MuI.result\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08951_ _01394_ _01401_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__nand2_1
XFILLER_170_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5115__A MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ _00483_ _00519_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__xnor2_1
XMuI._3988_ MuI._3039_ MuI._3054_ MuI._3059_ MuI._3087_ vssd1 vssd1 vccd1 vccd1 MuI._3088_
+ sky130_fd_sc_hd__and4bb_1
XMuI._6776_ MuI._2599_ MuI._2610_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2697_ sky130_fd_sc_hd__mux2_1
X_08882_ _06513_ _06611_ _04832_ _02420_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12820__A _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__A1 _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__A2 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5727_ MuI._1502_ MuI._1503_ MuI._1541_ MuI._1542_ vssd1 vssd1 vccd1 vccd1 MuI._1543_
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08733__B2 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ _00448_ _00449_ _00443_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a21o_1
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._607_ AuI.pe._145_ AuI.pe._022_ AuI.pe._041_ AuI.pe._142_ AuI.pe._159_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._160_ sky130_fd_sc_hd__a221o_1
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10978__C _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11436__A _04211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5658_ MuI._2860_ MuI._0246_ MuI._1005_ MuI._1004_ vssd1 vssd1 vccd1 vccd1 MuI._1467_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._5120__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _05627_ vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__clkbuf_4
XFILLER_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._538_ AuI.pe._095_ AuI.pe._370_ vssd1 vssd1 vccd1 vccd1 AuI.pe._096_ sky130_fd_sc_hd__nor2_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4609_ MuI._0311_ MuI._0303_ MuI._0309_ vssd1 vssd1 vccd1 vccd1 MuI._0313_ sky130_fd_sc_hd__nor3_1
X_09503_ _02112_ _02113_ _02114_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__o21ba_1
XMuI._5589_ MuI._1383_ MuI._1385_ MuI._1389_ vssd1 vssd1 vccd1 vccd1 MuI._1391_ sky130_fd_sc_hd__and3_1
X_06715_ _02356_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[4\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11155__B _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07695_ _00309_ _00312_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2b_1
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._469_ AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 AuI.pe._033_ sky130_fd_sc_hd__buf_2
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _02474_ _04165_ _00266_ _06564_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
XANTENNA__10843__A2 _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1396__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12045__A1 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13370__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _06663_ _04305_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__nand2_1
XFILLER_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5000__D MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ _03561_ _03928_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__nand2_2
XANTENNA_AuI._1409__B AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09296_ _01744_ _01806_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _00554_ _00558_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08178_ _00381_ _00388_ _00380_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07950__A2_N _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13098__A _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07129_ net127 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__buf_2
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__D _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _02815_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__and2_2
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08630__D _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10234__B _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__B1 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10071_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__buf_2
XANTENNA_AuI._1025__A0 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07543__B _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13481__B1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10973_ _03711_ _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__xnor2_4
XFILLER_189_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ _05134_ _02728_ _05584_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o21ai_1
XAuI._1050_ AuI._0110_ AuI._0248_ vssd1 vssd1 vccd1 vccd1 AuI._0261_ sky130_fd_sc_hd__xor2_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08077__D _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5695__A MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _05508_ _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nand2_1
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13233__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _05435_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor2_1
XFILLER_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10598__A1 AuI.result\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11525_ _04025_ _04149_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__a21oi_1
XFILLER_156_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3646__C MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._149_ FuI._012_ net155 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[20\] sky130_fd_sc_hd__dlxtn_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09486__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0903_ AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0123_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4866__A2_N MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11456_ _04232_ _04233_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nor2_1
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06903__A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4960_ MuI._0594_ MuI._0698_ vssd1 vssd1 vccd1 vccd1 MuI._0699_ sky130_fd_sc_hd__nor2_1
XFILLER_125_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07460__A1_N _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10407_ _00801_ _00802_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__and2b_1
XAuI._0834_ net107 vssd1 vssd1 vccd1 vccd1 AuI._0054_ sky130_fd_sc_hd__inv_2
X_11387_ _02566_ _02568_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__a21oi_1
XFILLER_180_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3911_ MuI._3008_ MuI._3010_ vssd1 vssd1 vccd1 vccd1 MuI._3011_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4891_ MuI._2754_ MuI._0228_ MuI._3371_ MuI._3000_ vssd1 vssd1 vccd1 vccd1 MuI._0623_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08219__A1_N _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08540__D _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ _03029_ _03027_ _03028_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nand3_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3842_ MuI._0867_ MuI._2787_ vssd1 vssd1 vccd1 vccd1 MuI._2942_ sky130_fd_sc_hd__nand2_1
XMuI._6630_ MuI._1766_ MuI._2535_ vssd1 vssd1 vccd1 vccd1 MuI._2536_ sky130_fd_sc_hd__nand2_1
XFILLER_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1016__A0 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05940_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI.pe._743__A2 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10269_ _00707_ _00708_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__or2_1
XFILLER_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6561_ MuI._2445_ MuI._2459_ vssd1 vssd1 vccd1 vccd1 MuI._2460_ sky130_fd_sc_hd__nand2_1
XFILLER_121_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3773_ MuI._2866_ vssd1 vssd1 vccd1 vccd1 MuI._2873_ sky130_fd_sc_hd__clkbuf_4
X_12008_ _04825_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5512_ MuI._3403_ MuI._3245_ MuI._3397_ MuI._0100_ vssd1 vssd1 vccd1 vccd1 MuI._1306_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1031__A3 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6492_ MuI._2380_ MuI._2383_ vssd1 vssd1 vccd1 vccd1 MuI._2384_ sky130_fd_sc_hd__nand2_1
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5443_ MuI._1217_ MuI._1227_ MuI._1166_ MuI._1228_ vssd1 vssd1 vccd1 vccd1 MuI._1231_
+ sky130_fd_sc_hd__a211o_1
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1317_ AuI._0276_ AuI._0307_ AuI._0294_ AuI._0389_ vssd1 vssd1 vccd1 vccd1 AuI._0514_
+ sky130_fd_sc_hd__a31o_1
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5374_ MuI._1101_ MuI._1103_ MuI._1102_ vssd1 vssd1 vccd1 vccd1 MuI._1155_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07480_ _00084_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__buf_4
XAuI._1248_ AuI._0438_ AuI._0313_ AuI._0421_ vssd1 vssd1 vccd1 vccd1 AuI._0450_ sky130_fd_sc_hd__o21a_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4325_ MuI._3255_ MuI._3280_ vssd1 vssd1 vccd1 vccd1 MuI._0002_ sky130_fd_sc_hd__nor2_1
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1179_ AuI._0266_ AuI._0384_ AuI._0269_ AuI._0267_ AuI._0176_ AuI._0206_ vssd1
+ vssd1 vccd1 vccd1 AuI._0385_ sky130_fd_sc_hd__mux4_1
XANTENNA_MuI._4613__B2 MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4256_ MuI._3227_ MuI._3228_ vssd1 vssd1 vccd1 vccd1 MuI._3356_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _01762_ _01764_ _01763_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08715__D _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10319__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _00714_ _00717_ _00718_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__nand3_1
XMuI._4187_ MuI._3215_ MuI._3254_ MuI._3286_ vssd1 vssd1 vccd1 vccd1 MuI._3287_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11250__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ _01344_ _01343_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__and2b_1
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08032_ _00646_ _00647_ _00648_ _00649_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__nand4_1
Xinput50 b_operand[21] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_6
Xinput61 b_operand[31] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_6
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6118__A1 MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3853__A MuI._2926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6118__B2 MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__B1 _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__A2_N _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09983_ _01304_ _01305_ _01306_ _01307_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__and4_1
XFILLER_131_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10054__B net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6828_ MuI._2700_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2746_ sky130_fd_sc_hd__and2b_1
X_08934_ _01497_ _01504_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nand2_1
XANTENNA__09843__B _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07509__A2 _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07644__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6759_ MuI._2676_ MuI._2677_ vssd1 vssd1 vccd1 vccd1 MuI._2678_ sky130_fd_sc_hd__nand2_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13365__B _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._474__C AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08865_ _01439_ _01440_ _01438_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__o21bai_1
XFILLER_96_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07816_ _00430_ _00432_ _00431_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a21o_1
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07363__B _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _01403_ _01404_ _01412_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__o21a_1
XANTENNA__09281__D _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._498__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07747_ _00360_ _00361_ _00363_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__or3_1
XFILLER_38_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3655__A2 MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07678_ _00286_ _00295_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ _02032_ _02034_ _02035_ _02036_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__o211a_1
XFILLER_13_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08906__C _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__B _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__B2 _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__B _00811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _06548_ _04509_ _00035_ _02291_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4959__A1_N MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__A2 _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _01789_ _01790_ _01793_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a21o_1
XANTENNA__11241__A2 _03828_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11310_ _00088_ _05187_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__nand2_1
XFILLER_193_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4907__A2 MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12290_ _05130_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06723__A _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ _03694_ _03828_ _04002_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5580__A2 MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5681__C MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3591__A1 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12741__A2 _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11172_ _00414_ _06622_ _05756_ _00785_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3913__D MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _04929_ _02916_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and2b_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A a_operand[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _02064_ net3 _02709_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__or3_2
XFILLER_0_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._489__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07704__D _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__A2 _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09122__A1 _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1102_ AuI._0225_ AuI._0227_ vssd1 vssd1 vccd1 vccd1 AuI._0312_ sky130_fd_sc_hd__nor2_1
XFILLER_204_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11804__A _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ _03556_ _03516_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__and2b_1
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1033_ AuI._0241_ AuI._0244_ AuI._0233_ vssd1 vssd1 vccd1 vccd1 AuI._0245_ sky130_fd_sc_hd__mux2_1
XANTENNA__07684__A1 _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07684__B2 _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4110_ MuI._3205_ MuI._3209_ vssd1 vssd1 vccd1 vccd1 MuI._3210_ sky130_fd_sc_hd__or2_1
XFILLER_92_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10887_ _03451_ _03453_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nand2_1
XMuI._5090_ MuI._0837_ MuI._0840_ MuI._0828_ MuI._0841_ vssd1 vssd1 vccd1 vccd1 MuI._0842_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _05289_ _05462_ _05463_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__nor3_2
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4041_ MuI._3133_ MuI._3134_ MuI._3139_ vssd1 vssd1 vccd1 vccd1 MuI._3141_ sky130_fd_sc_hd__a21o_1
XANTENNA__10139__B _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _05399_ _05287_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a21o_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4359__B1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11508_ _04287_ _04288_ _04269_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__a21o_1
XANTENNA__07729__A _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12980__A2 _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ _05340_ _05341_ _05343_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a21o_1
XFILLER_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5992_ MuI._1826_ MuI._1829_ MuI._1831_ MuI._1832_ MuI._1833_ vssd1 vssd1 vccd1
+ vccd1 MuI._1834_ sky130_fd_sc_hd__o311a_1
X_11439_ _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__or2b_1
XFILLER_172_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4943_ MuI._0576_ MuI._0679_ vssd1 vssd1 vccd1 vccd1 MuI._0681_ sky130_fd_sc_hd__nor2_1
XAuI._0817_ AuI._0036_ net13 vssd1 vssd1 vccd1 vccd1 AuI._0037_ sky130_fd_sc_hd__or2_1
XFILLER_125_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13109_ _05990_ _05991_ _05996_ _05997_ _06010_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__a221o_4
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4874_ MuI._0486_ MuI._0488_ vssd1 vssd1 vccd1 vccd1 MuI._0605_ sky130_fd_sc_hd__nor2_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ _05209_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__and3_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6613_ MuI._1645_ MuI._2516_ MuI._1460_ vssd1 vssd1 vccd1 vccd1 MuI._2518_ sky130_fd_sc_hd__mux2_1
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3825_ MuI._2906_ MuI._2923_ vssd1 vssd1 vccd1 vccd1 MuI._2925_ sky130_fd_sc_hd__and2b_1
XANTENNA__07464__A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__B1_N _04151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3885__A2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3756_ MuI._2055_ MuI._2852_ MuI.b_operand\[10\] MuI._2837_ vssd1 vssd1 vccd1
+ vccd1 MuI._2856_ sky130_fd_sc_hd__and4_1
XMuI._6544_ MuI._2439_ MuI._2432_ MuI._2438_ MuI._2441_ vssd1 vssd1 vccd1 vccd1 MuI._2442_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08650_ _01244_ _01243_ _01242_ _01228_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o211a_1
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._591__A AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07601_ _00217_ _00216_ _04843_ _04907_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__nand4_1
XFILLER_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3687_ MuI._2786_ vssd1 vssd1 vccd1 vccd1 MuI._2787_ sky130_fd_sc_hd__buf_2
XMuI._6475_ MuI._2364_ MuI._2365_ vssd1 vssd1 vccd1 vccd1 MuI._2366_ sky130_fd_sc_hd__or2_1
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08581_ _01182_ _01184_ _01196_ _01197_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__o211ai_4
XFILLER_81_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5426_ MuI._1206_ MuI._1211_ vssd1 vssd1 vccd1 vccd1 MuI._1212_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12799__A2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ net116 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__buf_4
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07911__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__A _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5357_ MuI._1129_ MuI._1130_ MuI._1135_ vssd1 vssd1 vccd1 vccd1 MuI._1136_ sky130_fd_sc_hd__a21o_1
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08726__C net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11433__B _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ net117 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__clkbuf_4
XMuI._4308_ MuI._3395_ MuI._3406_ MuI._3407_ vssd1 vssd1 vccd1 vccd1 MuI._3408_ sky130_fd_sc_hd__a21bo_1
XFILLER_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09202_ _01817_ _01818_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__o21bai_1
XMuI._5288_ MuI._0992_ MuI._1059_ vssd1 vssd1 vccd1 vccd1 MuI._1060_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _06598_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__buf_6
XMuI._4239_ MuI._3233_ MuI._3234_ MuI._3252_ vssd1 vssd1 vccd1 vccd1 MuI._3339_ sky130_fd_sc_hd__o21a_1
XFILLER_176_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ _01727_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__inv_2
XFILLER_148_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _02334_ _00032_ _06611_ _01332_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__a22o_1
XANTENNA__07639__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08461__C _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _00629_ _00631_ _00632_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a21bo_1
XFILLER_163_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10065__A _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._766__A AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ _02041_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__and2_1
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4522__B1 MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _01486_ _01491_ _01485_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a21bo_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _02555_ _02541_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__xnor2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5303__A MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10498__B1 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _01462_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xnor2_1
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ net120 net44 _00271_ _04229_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__and4_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _03395_ _03398_ _03396_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o21bai_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6027__B1 MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _04591_ _04592_ _04420_ _04422_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__a211o_1
XANTENNA__06718__A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A2 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11998__B1 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _03460_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__a21o_1
XFILLER_201_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13460_ _01330_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
XFILLER_201_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10672_ _03386_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21o_1
XFILLER_167_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _02795_ _05249_ _05017_ _05260_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__o31ai_1
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _06304_ _02699_ _01322_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__o21ai_4
XFILLER_182_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11997__C _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08652__B _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ _03389_ _03454_ _05391_ _06546_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__nand4_1
XFILLER_166_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3493__A MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5553__A2 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _05077_ _05111_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nor3_4
XFILLER_154_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12714__A2 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _03754_ _03947_ _03983_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a211oi_4
XAuI._1651_ AuI._0603_ AuI._0692_ AuI.operand_a\[26\] AuI._0258_ vssd1 vssd1 vccd1
+ vccd1 AuI._0006_ sky130_fd_sc_hd__a211o_1
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12902__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12190__A3 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _02539_ _05959_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__nand2_1
XAuI._1582_ AuI._0755_ AuI._0756_ vssd1 vssd1 vccd1 vccd1 AuI._0757_ sky130_fd_sc_hd__nor2_1
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10106_ _05467_ _03346_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__or2b_1
XANTENNA__07284__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3940__B MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11086_ _02530_ _02544_ _02564_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__nor3_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3610_ MuI._2055_ vssd1 vssd1 vccd1 vccd1 MuI._2066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_103_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08099__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4590_ MuI._1296_ MuI._1791_ MuI._3362_ MuI._2829_ vssd1 vssd1 vccd1 vccd1 MuI._0292_
+ sky130_fd_sc_hd__and4_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10037_ _02064_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__nor2_2
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3541_ MuI._1296_ vssd1 vssd1 vccd1 vccd1 MuI._1307_ sky130_fd_sc_hd__buf_2
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6743__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6260_ MuI._0570_ MuI._1318_ MuI._1813_ MuI._0339_ vssd1 vssd1 vccd1 vccd1 MuI._2129_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3472_ MuI._0471_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._0548_ sky130_fd_sc_hd__nand2_1
XFILLER_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5211_ MuI._0969_ MuI._0972_ MuI._0973_ MuI._0974_ vssd1 vssd1 vccd1 vccd1 MuI._0975_
+ sky130_fd_sc_hd__a211o_1
X_11988_ _04804_ _04805_ _04770_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__o21a_1
XFILLER_205_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__A2 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6191_ MuI._2051_ MuI._2052_ MuI._0867_ MuI._2627_ vssd1 vssd1 vccd1 vccd1 MuI._2053_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA_MuI._3668__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ MuI.result\[4\] _02736_ _02707_ _02764_ _03676_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5586__C MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5142_ MuI._2875_ MuI._2341_ MuI._0085_ MuI._2873_ vssd1 vssd1 vccd1 vccd1 MuI._0899_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1016_ net67 net35 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0228_ sky130_fd_sc_hd__mux2_1
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08265__D _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5073_ MuI._0819_ MuI._0822_ vssd1 vssd1 vccd1 vccd1 MuI._0824_ sky130_fd_sc_hd__xor2_1
XFILLER_192_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _05335_ _05398_ _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12402__A1 _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__B _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4024_ MuI._3121_ MuI._3122_ MuI._3085_ MuI._3086_ vssd1 vssd1 vccd1 vccd1 MuI._3124_
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07459__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5544__A2 MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09096__D net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5975_ MuI._1809_ MuI._1815_ vssd1 vssd1 vccd1 vccd1 MuI._1816_ sky130_fd_sc_hd__nand2_1
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5107__B MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3553__D MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4926_ MuI._0452_ MuI._0661_ vssd1 vssd1 vccd1 vccd1 MuI._0662_ sky130_fd_sc_hd__xor2_2
XFILLER_141_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _02451_ _02452_ _02466_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11709__A _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._786_ AuI.pe._323_ AuI.pe._324_ AuI.pe._325_ AuI.pe._319_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._327_ sky130_fd_sc_hd__o31ai_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07194__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4857_ MuI._0517_ MuI._0518_ MuI._0519_ vssd1 vssd1 vccd1 vccd1 MuI._0586_ sky130_fd_sc_hd__a21oi_1
X_09751_ _02322_ _02395_ _02397_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__nor3_1
XFILLER_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06963_ _05025_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__buf_6
XANTENNA__10332__B _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3808_ MuI._1010_ MuI._1472_ MuI._2836_ MuI._2838_ vssd1 vssd1 vccd1 vccd1 MuI._2908_
+ sky130_fd_sc_hd__and4_1
X_08702_ _01200_ _01201_ _01319_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__nand3_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4788_ MuI._0507_ MuI._0509_ vssd1 vssd1 vccd1 vccd1 MuI._0510_ sky130_fd_sc_hd__and2b_1
XANTENNA_AuI.pe._570__B1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ _02219_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__or2_1
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06894_ net123 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__buf_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6527_ MuI._2422_ vssd1 vssd1 vccd1 vccd1 MuI._2423_ sky130_fd_sc_hd__inv_2
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3739_ MuI._1461_ MuI._2055_ MuI._2836_ MuI._2838_ vssd1 vssd1 vccd1 vccd1 MuI._2839_
+ sky130_fd_sc_hd__and4_1
X_08633_ _01250_ _01081_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__xnor2_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6458_ MuI._2343_ MuI._2345_ vssd1 vssd1 vccd1 vccd1 MuI._2347_ sky130_fd_sc_hd__xor2_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09098__B1 _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08564_ _01129_ _01131_ _01181_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__o21a_1
XFILLER_82_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5409_ MuI._1134_ MuI._1133_ MuI._1132_ vssd1 vssd1 vccd1 vccd1 MuI._1193_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12259__B _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ net118 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__buf_4
XMuI._6389_ MuI._1966_ MuI._1969_ vssd1 vssd1 vccd1 vccd1 MuI._2271_ sky130_fd_sc_hd__or2_1
XANTENNA__08845__B1 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ _01108_ _01109_ _01111_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__nor3_1
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07446_ _00062_ _00040_ _06612_ _00063_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__a22oi_1
XFILLER_210_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07377_ _06619_ _06627_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and2b_1
XFILLER_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ _01612_ _01611_ _01613_ _01614_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__or4b_2
XFILLER_164_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1417__B AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _01566_ _01590_ _01663_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__o211a_2
XANTENNA__12425__D _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08306__B1_N _00923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10523__A _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09949_ _02341_ _02340_ _02610_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a31o_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13121__A2 _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ FuI.Integer\[21\] _04627_ _02731_ AuI.result\[21\] vssd1 vssd1 vccd1 vccd1
+ _05851_ sky130_fd_sc_hd__a22o_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09876__A2 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ _04527_ _04529_ _04528_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__o21bai_1
XFILLER_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12891_ _05744_ _05742_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or2b_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ AuI.result\[11\] _02732_ _04648_ _02935_ vssd1 vssd1 vccd1 vccd1 _04650_
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5471__A1 MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _00281_ _03443_ _05036_ _00534_ vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__nand4_2
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10643__B1 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ _03442_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__nor2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08663__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13443_ _06355_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__xnor2_1
X_10655_ _03368_ _03369_ _03165_ _03169_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o211ai_1
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07279__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _06276_ _06285_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__or2_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10586_ _03294_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nand2_1
XFILLER_182_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12325_ _05059_ _05061_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4734__B1 MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12256_ _02980_ _03047_ _06477_ _00281_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a22o_1
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5760_ MuI._1576_ MuI._1577_ MuI._1575_ vssd1 vssd1 vccd1 vccd1 MuI._1579_ sky130_fd_sc_hd__a21bo_1
X_11207_ _03964_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_1
XAuI._1634_ AuI._0693_ AuI._0795_ AuI._0798_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0799_
+ sky130_fd_sc_hd__o22a_1
X_12187_ _02795_ _05018_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__nand2_1
XAuI.pe._640_ AuI.pe.significand\[12\] AuI.pe._004_ AuI.pe._022_ AuI.pe._170_ AuI.pe._190_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._191_ sky130_fd_sc_hd__a221o_1
XFILLER_110_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4711_ MuI._0423_ MuI._0424_ MuI.b_operand\[14\] MuI._3363_ vssd1 vssd1 vccd1
+ vccd1 MuI._0425_ sky130_fd_sc_hd__and4bb_1
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3670__B MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5691_ MuI._1500_ MuI._1501_ MuI._1480_ MuI._1481_ vssd1 vssd1 vccd1 vccd1 MuI._1503_
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11138_ _03888_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a21o_1
XAuI._1565_ AuI._0701_ AuI._0738_ AuI._0742_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0743_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_MuI._6039__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._571_ AuI.pe._106_ AuI.pe._023_ AuI.pe._042_ AuI.pe._102_ AuI.pe._126_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._127_ sky130_fd_sc_hd__a221o_1
XANTENNA_MuI._4485__C MuI._0175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4642_ MuI._0342_ MuI._0346_ MuI._0348_ vssd1 vssd1 vccd1 vccd1 MuI._0349_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11069_ _03814_ _03815_ _03639_ _03641_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__a211o_1
XFILLER_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1496_ AuI._0564_ AuI._0566_ vssd1 vssd1 vccd1 vccd1 AuI._0682_ sky130_fd_sc_hd__and2_1
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12320__B1 _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4573_ MuI._0264_ MuI._0265_ vssd1 vssd1 vccd1 vccd1 MuI._0274_ sky130_fd_sc_hd__and2b_1
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4782__A MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6312_ MuI._2161_ MuI._2162_ MuI._2184_ vssd1 vssd1 vccd1 vccd1 MuI._2186_ sky130_fd_sc_hd__or3_1
XFILLER_92_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3524_ MuI._0350_ MuI._0889_ MuI._0746_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._1120_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4713__A1_N MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6243_ MuI._1153_ MuI._1032_ MuI._1483_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._2111_
+ sky130_fd_sc_hd__a22oi_1
XMuI._3455_ MuI.b_operand\[22\] vssd1 vssd1 vccd1 vccd1 MuI._0361_ sky130_fd_sc_hd__clkbuf_2
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11426__A2 _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__C net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ net41 vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6174_ MuI.a_operand\[19\] MuI._1461_ MuI._1296_ MuI.b_operand\[15\] vssd1 vssd1
+ vccd1 vccd1 MuI._2035_ sky130_fd_sc_hd__and4_1
X_08280_ _00580_ _00581_ _00583_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__o21a_1
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5125_ MuI._0871_ MuI._0879_ MuI._0880_ vssd1 vssd1 vccd1 vccd1 MuI._0881_ sky130_fd_sc_hd__nand3_1
X_07231_ _06523_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5056_ MuI._0800_ MuI._0804_ vssd1 vssd1 vccd1 vccd1 MuI._0805_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07189__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07162_ net116 vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__buf_6
XMuI._4007_ MuI._3105_ MuI._3106_ vssd1 vssd1 vccd1 vccd1 MuI._3107_ sky130_fd_sc_hd__nor2_1
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07093_ _04994_ _06284_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__and2_1
XFILLER_118_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6190__A2 MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06821__A _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3861__A MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5958_ MuI._0730_ MuI._1777_ MuI._1779_ vssd1 vssd1 vccd1 vccd1 MuI._1797_ sky130_fd_sc_hd__or3_1
XANTENNA__13351__A2 _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4909_ MuI._0640_ MuI._0642_ vssd1 vssd1 vccd1 vccd1 MuI._0643_ sky130_fd_sc_hd__nor2_1
X_09803_ net110 net109 net132 net127 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__and4_1
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5889_ MuI._1654_ MuI._1657_ vssd1 vssd1 vccd1 vccd1 MuI._1721_ sky130_fd_sc_hd__or2b_1
XANTENNA__11158__B _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12969__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _00298_ _00316_ _00315_ _00308_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a211o_1
XAuI.pe._769_ AuI.pe._056_ AuI.pe._225_ AuI.pe._296_ AuI.pe._303_ AuI.pe._312_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._313_ sky130_fd_sc_hd__a2111o_1
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ _02378_ _02379_ _02604_ _03917_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__o211a_1
XANTENNA__13103__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06946_ _04843_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07688__A2_N _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07652__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09665_ _02289_ _02290_ _02303_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a21o_1
XANTENNA__07869__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _04100_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__clkbuf_4
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07869__B2 _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ _01025_ _01024_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__and2b_1
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08530__A2 _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__B1 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09596_ _02228_ _02230_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__o21ba_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _03335_ _03884_ _01145_ _01148_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a22oi_1
XFILLER_196_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3739__C MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11902__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08294__A1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _01094_ _01095_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__xnor2_2
XANTENNA__08294__B2 _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07429_ _04574_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__buf_4
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__A _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _03005_ _03042_ _03040_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__o21ai_2
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__A1 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _03063_ _03064_ _00762_ _00764_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__o211a_1
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4716__B1 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _04906_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__xor2_1
XFILLER_151_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07827__A _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _05988_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__nand2_1
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06731__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3771__A MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09546__A1 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09546__B2 _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _04751_ _04753_ _04862_ _04863_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__o211ai_4
XFILLER_105_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4586__B MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07265__C _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1350_ AuI._0543_ AuI._0544_ vssd1 vssd1 vccd1 vccd1 AuI._0545_ sky130_fd_sc_hd__and2b_1
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _05829_ _05830_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__nand2_1
XAuI._1281_ AuI._0455_ AuI._0468_ vssd1 vssd1 vccd1 vccd1 AuI._0481_ sky130_fd_sc_hd__nand2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__A2 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07281__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _02856_ _02868_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__nor2_1
XANTENNA__08808__D _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _03489_ _04625_ _04631_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a21o_1
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output102_A net102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _00678_ _06603_ _06605_ _03539_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a22o_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06906__A _04413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__B _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _00000_ _06682_ _05574_ _03425_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__nand4_1
XFILLER_187_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11687_ _04360_ _04304_ _04482_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a211o_1
XFILLER_128_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13426_ _06334_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__xnor2_1
X_10638_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__nor2_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13357_ _02751_ _06221_ _06223_ _06257_ _06269_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__a311o_4
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ _03276_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0996_ AuI._0100_ AuI._0207_ vssd1 vssd1 vccd1 vccd1 AuI._0208_ sky130_fd_sc_hd__xnor2_4
XFILLER_170_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0896__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6861_ MuI._2762_ MuI._2763_ vssd1 vssd1 vccd1 vccd1 MuI._2764_ sky130_fd_sc_hd__xnor2_1
X_12308_ _03013_ _05959_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__nand2_1
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13288_ _06197_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__inv_2
XMuI._5812_ MuI._1633_ MuI._1634_ MuI._1545_ MuI._1547_ vssd1 vssd1 vccd1 vccd1 MuI._1636_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6792_ MuI._2707_ MuI._2711_ MuI._2712_ MuI._2713_ vssd1 vssd1 vccd1 vccd1 MuI._2714_
+ sky130_fd_sc_hd__and4b_1
X_12239_ _04936_ _04935_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or2b_1
XANTENNA__10163__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5743_ MuI._3000_ MuI._2754_ MuI._0110_ MuI.a_operand\[1\] vssd1 vssd1 vccd1
+ vccd1 MuI._1561_ sky130_fd_sc_hd__and4_1
XAuI._1617_ AuI.pe.Significand\[17\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0786_
+ sky130_fd_sc_hd__or2_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._623_ AuI.pe._046_ AuI.pe._133_ AuI.pe._173_ AuI.pe._030_ AuI.pe._174_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._175_ sky130_fd_sc_hd__a221o_1
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06800_ _03271_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__buf_4
XMuI._5674_ MuI._2853_ MuI._2854_ MuI.a_operand\[7\] MuI.a_operand\[6\] vssd1 vssd1
+ vccd1 vccd1 MuI._1485_ sky130_fd_sc_hd__and4_1
XFILLER_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1548_ AuI._0701_ AuI._0724_ AuI._0728_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0729_
+ sky130_fd_sc_hd__o22a_1
X_07780_ _06466_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__buf_4
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._554_ AuI.pe._055_ AuI.pe._086_ AuI.pe._110_ vssd1 vssd1 vccd1 vccd1 AuI.pe._111_
+ sky130_fd_sc_hd__a21o_1
XMuI._4625_ MuI._0329_ MuI._0330_ MuI.b_operand\[11\] MuI._2790_ vssd1 vssd1 vccd1
+ vccd1 MuI._0331_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07472__A _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 Operation[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
X_06731_ _02528_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__buf_6
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1479_ AuI._0422_ AuI._0424_ AuI._0428_ vssd1 vssd1 vccd1 vccd1 AuI._0665_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10610__B _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._485_ AuI.pe.significand\[1\] AuI.pe.significand\[0\] AuI.pe.significand\[2\]
+ AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 AuI.pe._048_ sky130_fd_sc_hd__or4_1
XMuI._4556_ MuI._0176_ MuI._0197_ MuI._0199_ vssd1 vssd1 vccd1 vccd1 MuI._0255_ sky130_fd_sc_hd__a21o_1
X_09450_ _02068_ _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3507_ MuI._0911_ MuI._0922_ vssd1 vssd1 vccd1 vccd1 MuI._0933_ sky130_fd_sc_hd__nand2_1
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08401_ _02593_ _02658_ _04778_ _06603_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__and4_1
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4487_ MuI._0172_ MuI._0178_ vssd1 vssd1 vccd1 vccd1 MuI._0179_ sky130_fd_sc_hd__xnor2_1
X_09381_ _01997_ _01998_ net122 _04035_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and4bb_1
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6226_ MuI._2086_ MuI._2091_ vssd1 vssd1 vccd1 vccd1 MuI._2092_ sky130_fd_sc_hd__xnor2_1
XMuI._3438_ MuI._0108_ MuI._0152_ MuI._0163_ vssd1 vssd1 vccd1 vccd1 MuI._0174_ sky130_fd_sc_hd__a21bo_1
X_08332_ _00947_ _00948_ _00949_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__nor3_1
XFILLER_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09473__B1 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06816__A _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6157_ MuI._2014_ MuI._2015_ vssd1 vssd1 vccd1 vccd1 MuI._2016_ sky130_fd_sc_hd__nor2_1
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08263_ _00571_ _00573_ _00572_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__o21ai_1
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout133_A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5108_ MuI._0860_ MuI._0861_ vssd1 vssd1 vccd1 vccd1 MuI._0862_ sky130_fd_sc_hd__nor2_1
XFILLER_165_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4946__B1 MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ net66 vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__clkbuf_4
XMuI._6088_ MuI._1927_ MuI._1928_ MuI._1938_ vssd1 vssd1 vccd1 vccd1 MuI._1940_ sky130_fd_sc_hd__nand3_1
XFILLER_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08453__D _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ _00810_ _00811_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__xor2_2
XFILLER_193_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5039_ MuI._0418_ MuI._0547_ MuI._0551_ MuI._0784_ MuI._0785_ vssd1 vssd1 vccd1
+ vccd1 MuI._0786_ sky130_fd_sc_hd__a221o_1
XANTENNA__09776__A1 _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B2 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ net127 vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__buf_4
XFILLER_106_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07076_ _04467_ _06067_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11169__A _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13324__A2 _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07366__B _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3921__A1 MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__B1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11335__B2 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3921__B2 MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08200__A1 _00664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _00593_ _00594_ _00595_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__or3_2
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10801__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07382__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _02359_ _02360_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11616__B _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06929_ _04660_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _02284_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__nor2_1
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08628__D _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _02209_ _02210_ _02204_ _02208_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__o211a_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._810__D_N AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08939__A2_N _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11610_ _01146_ _00002_ _06561_ _01147_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a22oi_1
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12063__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12590_ _05451_ _05452_ _05444_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__a21o_1
XANTENNA__08267__B2 _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09464__B1 _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06726__A _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _02773_ _04163_ _01891_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__o21a_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__B1 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _04248_ _04249_ _04184_ _04185_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__o211ai_4
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._096_ FuI._037_ net104 FuI._056_ vssd1 vssd1 vccd1 vccd1 FuI._057_ sky130_fd_sc_hd__and3_1
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13211_ _06116_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__nand2_1
XFILLER_171_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09767__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _03118_ _03120_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__nand2_1
XAuI._0850_ net8 vssd1 vssd1 vccd1 vccd1 AuI._0070_ sky130_fd_sc_hd__inv_2
XFILLER_164_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07557__A net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ _06041_ _06044_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input63_A b_operand[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _00877_ _00878_ _06561_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__and4_1
XFILLER_124_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13073_ _03809_ _05520_ _05969_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21o_1
XFILLER_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10285_ _02960_ _02961_ _02972_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__and3_1
XFILLER_152_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12024_ _04842_ _04844_ _04831_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11877__A2 _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1402_ AuI._0579_ AuI._0591_ vssd1 vssd1 vccd1 vccd1 AuI._0592_ sky130_fd_sc_hd__nand2_1
XANTENNA__08742__A2 _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._507__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11807__A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07292__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1333_ AuI._0507_ AuI._0508_ AuI._0520_ AuI._0521_ vssd1 vssd1 vccd1 vccd1 AuI._0529_
+ sky130_fd_sc_hd__or4_1
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4410_ MuI._0084_ MuI._0092_ MuI._0093_ vssd1 vssd1 vccd1 vccd1 MuI._0094_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5221__A MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5390_ MuI._1119_ MuI._1171_ vssd1 vssd1 vccd1 vccd1 MuI._1172_ sky130_fd_sc_hd__or2_1
XFILLER_207_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1264_ AuI._0442_ AuI._0451_ AuI._0463_ vssd1 vssd1 vccd1 vccd1 AuI._0465_ sky130_fd_sc_hd__and3_1
XFILLER_19_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _05721_ _05720_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__or2b_1
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4341_ MuI.a_operand\[22\] MuI._0559_ MuI._0017_ MuI._0018_ vssd1 vssd1 vccd1
+ vccd1 MuI._0019_ sky130_fd_sc_hd__and4_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1195_ AuI._0256_ AuI._0377_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0401_ sky130_fd_sc_hd__and3_1
X_12857_ _05655_ _05658_ _05739_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__or3_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12638__A _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4272_ MuI._3371_ vssd1 vssd1 vccd1 vccd1 MuI._3372_ sky130_fd_sc_hd__buf_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08258__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ _04612_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__xnor2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08258__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12788_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
XMuI._6011_ MuI._1813_ MuI._2066_ MuI._2916_ MuI._1318_ vssd1 vssd1 vccd1 vccd1 MuI._1855_
+ sky130_fd_sc_hd__a22oi_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__B _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _04406_ _04408_ _04407_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o21bai_1
XANTENNA_MuI._6393__A2 MuI._1975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07481__A2 _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13409_ _03842_ _05917_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__nand2_1
XFILLER_143_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07467__A _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._0979_ AuI._0165_ AuI._0167_ AuI._0117_ vssd1 vssd1 vccd1 vccd1 AuI._0191_ sky130_fd_sc_hd__a21oi_2
XFILLER_131_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__B _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6844_ MuI._2694_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2755_ sky130_fd_sc_hd__and2b_1
X_08950_ _01395_ _01400_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__or2b_1
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07901_ _00501_ _00518_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__xnor2_4
XMuI._6775_ MuI._2632_ MuI._2636_ MuI._2641_ vssd1 vssd1 vccd1 vccd1 MuI._2696_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3987_ MuI._3046_ MuI._3047_ MuI._3052_ vssd1 vssd1 vccd1 vccd1 MuI._3087_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._5115__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08881_ _06519_ _06515_ _04767_ net10 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__and4_1
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12820__B _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5726_ MuI._1539_ MuI._1540_ MuI._1048_ MuI._1504_ vssd1 vssd1 vccd1 vccd1 MuI._1542_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08733__A2 _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__A _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _00443_ _00448_ _00449_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__nand3_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07914__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._606_ AuI.pe._158_ AuI.pe._025_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._159_
+ sky130_fd_sc_hd__a21o_1
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08298__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5657_ MuI._1009_ MuI._1011_ MuI._1013_ vssd1 vssd1 vccd1 vccd1 MuI._1466_ sky130_fd_sc_hd__nand3_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__D _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _00377_ _00379_ _00378_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__a21o_1
XFILLER_84_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._537_ AuI.pe.significand\[15\] vssd1 vssd1 vccd1 vccd1 AuI.pe._095_ sky130_fd_sc_hd__inv_2
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4608_ MuI._0303_ MuI._0309_ MuI._0311_ vssd1 vssd1 vccd1 vccd1 MuI._0312_ sky130_fd_sc_hd__o21a_1
X_09502_ _02539_ _04186_ _02049_ _02048_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._5131__A MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06714_ _02345_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__and3_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5588_ MuI._1383_ MuI._1385_ MuI._1389_ vssd1 vssd1 vccd1 vccd1 MuI._1390_ sky130_fd_sc_hd__a21o_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07694_ _00309_ _00310_ _00311_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__or3_1
XFILLER_198_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._468_ AuI.pe._020_ AuI.pe._023_ AuI.pe._027_ AuI.pe._029_ AuI.pe._032_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe.Significand\[1\] sky130_fd_sc_hd__a221o_1
XFILLER_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4539_ MuI._0230_ MuI._0233_ MuI._0235_ vssd1 vssd1 vccd1 vccd1 MuI._0236_ sky130_fd_sc_hd__o21a_1
X_09433_ _06520_ _06513_ _00271_ _04229_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__nand4_1
XFILLER_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4970__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _01966_ _01969_ _01967_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__o21ba_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4092__B1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12045__A2 _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6209_ MuI._2063_ MuI._2071_ MuI._2072_ vssd1 vssd1 vccd1 vccd1 MuI._2073_ sky130_fd_sc_hd__nand3_1
XFILLER_33_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08315_ _00909_ _00932_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__or2_1
X_09295_ _01898_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__nand2_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08246_ _00843_ _00839_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__or2b_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _00788_ _00794_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11556__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07128_ net60 vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13098__B _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4848__C MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07059_ _06056_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11308__A1 _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__B2 _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__buf_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1025__A1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07543__C _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ _00502_ _04316_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nand2_1
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _02129_ _02854_ _02855_ _04011_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__o211ai_1
XANTENNA__11492__B1 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11362__A _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _05416_ _05507_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5695__B MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3496__A MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ _05423_ _05424_ _05433_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and3_1
XFILLER_200_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10598__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__B1 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11524_ _04148_ _04147_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__and2b_2
XFILLER_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3646__D MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFuI._148_ FuI._011_ net154 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[19\] sky130_fd_sc_hd__dlxtn_1
XAuI._0902_ AuI._0121_ vssd1 vssd1 vccd1 vccd1 AuI._0122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09486__B _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ _06606_ _06601_ _06537_ _00385_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__and4_1
XFILLER_172_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11547__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFuI._079_ FuI.a_operand\[26\] FuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 FuI._044_
+ sky130_fd_sc_hd__nor2_1
XFILLER_137_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10406_ _03043_ _03103_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__xor2_2
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0833_ net66 vssd1 vssd1 vccd1 vccd1 AuI._0053_ sky130_fd_sc_hd__inv_2
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3910_ MuI._2927_ MuI._2934_ MuI._3009_ vssd1 vssd1 vccd1 vccd1 MuI._3010_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4138__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4138__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _03744_ _05660_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nand2_1
XMuI._4890_ MuI._1296_ MuI._1791_ MuI._3245_ MuI._0304_ vssd1 vssd1 vccd1 vccd1 MuI._0622_
+ sky130_fd_sc_hd__and4_1
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _03027_ _03028_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4120__A MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3841_ MuI._2938_ MuI._2940_ vssd1 vssd1 vccd1 vccd1 MuI._2941_ sky130_fd_sc_hd__nor2_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _05950_ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI._1016__A1 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10268_ _00707_ _00708_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
XFILLER_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6560_ MuI._2457_ MuI._2458_ vssd1 vssd1 vccd1 vccd1 MuI._2459_ sky130_fd_sc_hd__nor2_1
X_12007_ _04713_ _04715_ _04826_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a21oi_1
XMuI._3772_ MuI._1483_ MuI._2871_ vssd1 vssd1 vccd1 vccd1 MuI._2872_ sky130_fd_sc_hd__nand2_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _02216_ _03993_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__or2b_1
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5511_ MuI._3268_ MuI._3371_ vssd1 vssd1 vccd1 vccd1 MuI._1305_ sky130_fd_sc_hd__nand2_1
XFILLER_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6491_ MuI._2381_ MuI._2382_ vssd1 vssd1 vccd1 vccd1 MuI._2383_ sky130_fd_sc_hd__xor2_1
XANTENNA__10160__B _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6047__A MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5442_ MuI._1217_ MuI._1227_ MuI._1166_ MuI._1228_ vssd1 vssd1 vccd1 vccd1 MuI._1229_
+ sky130_fd_sc_hd__a211oi_2
XAuI._1316_ AuI._0508_ AuI._0512_ AuI._0507_ vssd1 vssd1 vccd1 vccd1 AuI._0513_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08846__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5373_ MuI._1101_ MuI._1102_ MuI._1103_ vssd1 vssd1 vccd1 vccd1 MuI._1154_ sky130_fd_sc_hd__and3_1
X_12909_ _05699_ _05703_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XAuI._1247_ AuI._0306_ AuI._0308_ vssd1 vssd1 vccd1 vccd1 AuI._0449_ sky130_fd_sc_hd__and2_1
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4324_ MuI._3255_ MuI._3280_ vssd1 vssd1 vccd1 vccd1 MuI._0001_ sky130_fd_sc_hd__and2_1
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11272__A _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09428__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1178_ AuI._0199_ AuI._0200_ AuI._0226_ vssd1 vssd1 vccd1 vccd1 AuI._0384_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4613__A2 MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4255_ MuI._3353_ MuI._3354_ vssd1 vssd1 vccd1 vccd1 MuI._3355_ sky130_fd_sc_hd__nand2_1
XFILLER_203_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _00444_ _00550_ _00715_ _00716_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__a22o_1
XMuI._4186_ MuI._2834_ MuI._3212_ MuI._3213_ vssd1 vssd1 vccd1 vccd1 MuI._3286_ sky130_fd_sc_hd__and3_1
XFILLER_175_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__C _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09080_ _02528_ _00085_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__nand2_1
XFILLER_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4014__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08031_ _00564_ _00585_ _00579_ _00584_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__o211ai_2
XFILLER_175_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 b_operand[12] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_6
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 b_operand[22] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_4
Xinput62 b_operand[3] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_4
XFILLER_156_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6118__A2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08403__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ _01304_ _01305_ _01306_ _01307_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22oi_4
XFILLER_171_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6827_ MuI._2745_ vssd1 vssd1 vccd1 vccd1 MuI.result\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08933_ _01501_ _01498_ _01502_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__or3_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6758_ MuI._2643_ MuI._2647_ MuI._2675_ vssd1 vssd1 vccd1 vccd1 MuI._2677_ sky130_fd_sc_hd__a21o_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08864_ _01283_ _01281_ _01282_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__or3_1
XANTENNA__10351__A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5709_ MuI._2484_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._1523_ sky130_fd_sc_hd__nand2_1
XFILLER_111_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07815_ _00430_ _00431_ _00432_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__nand3_1
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6689_ MuI._2600_ vssd1 vssd1 vccd1 vccd1 MuI._2601_ sky130_fd_sc_hd__inv_2
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _01403_ _01404_ _01412_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nor3_4
XFILLER_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4301__A1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07746_ _00360_ _00361_ _00363_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08756__A _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07660__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _00293_ _00294_ vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__nor2_1
XFILLER_198_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _01957_ _01956_ _01924_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13215__A1 _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__D _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07693__A2 _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _01936_ _01928_ _01935_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__nand3_1
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _01889_ _01894_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a21o_1
XFILLER_194_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08229_ _00635_ _00636_ _00637_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__a21oi_2
XFILLER_181_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06723__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _03827_ _03824_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__and2b_2
XFILLER_181_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5681__D MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13350__A1_N _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3591__A2 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _02658_ _00385_ _00783_ _02593_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a22oi_2
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ _02796_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__inv_2
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _02118_ _03928_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__o21a_1
XFILLER_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input26_A a_operand[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._489__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1101_ AuI._0272_ AuI._0270_ AuI._0175_ vssd1 vssd1 vccd1 vccd1 AuI._0311_ sky130_fd_sc_hd__mux2_1
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09122__A2 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ _03820_ _04262_ _03532_ _03530_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__a31o_1
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1032_ AuI._0242_ AuI._0243_ AuI._0205_ vssd1 vssd1 vccd1 vccd1 AuI._0244_ sky130_fd_sc_hd__mux2_1
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _03617_ _03618_ _03598_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a21o_1
XANTENNA__07684__A2 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _03831_ _05134_ _05437_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and3_1
XFILLER_169_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4040_ MuI._3133_ MuI._3134_ MuI._3139_ vssd1 vssd1 vccd1 vccd1 MuI._3140_ sky130_fd_sc_hd__nand3_1
XFILLER_185_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13303__A1_N _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_8 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__A _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12965__B1 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06914__A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4359__A1 MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4359__B2 MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _04269_ _04287_ _04288_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nand3_1
XFILLER_172_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07729__B _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ _05340_ _05341_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__nand3_1
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output94_A net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5991_ MuI._1817_ MuI._1825_ vssd1 vssd1 vccd1 vccd1 MuI._1833_ sky130_fd_sc_hd__or2_1
X_11438_ _04212_ _04213_ _04076_ _04207_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a211o_1
XFILLER_99_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4942_ MuI._2484_ MuI._0168_ MuI._0574_ MuI._0575_ vssd1 vssd1 vccd1 vccd1 MuI._0679_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_113_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0816_ net119 vssd1 vssd1 vccd1 vccd1 AuI._0036_ sky130_fd_sc_hd__inv_2
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11369_ _04094_ _04095_ _04138_ _04139_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__a22oi_4
XFILLER_180_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4873_ MuI._0577_ MuI._0583_ vssd1 vssd1 vccd1 vccd1 MuI._0604_ sky130_fd_sc_hd__or2b_1
X_13108_ _03315_ _05999_ _06000_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__a31o_1
XFILLER_113_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6612_ MuI._1642_ MuI._1643_ MuI._2515_ vssd1 vssd1 vccd1 vccd1 MuI._2516_ sky130_fd_sc_hd__o21ba_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3824_ MuI._2906_ MuI._2923_ vssd1 vssd1 vccd1 vccd1 MuI._2924_ sky130_fd_sc_hd__xnor2_2
XFILLER_112_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11267__A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _03489_ _05929_ _05930_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__a31o_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13185__C _06091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6543_ MuI._2414_ MuI._2427_ MuI._2437_ vssd1 vssd1 vccd1 vccd1 MuI._2441_ sky130_fd_sc_hd__o21bai_1
XMuI._3755_ MuI._2852_ MuI._2853_ MuI._2854_ MuI._2055_ vssd1 vssd1 vccd1 vccd1 MuI._2855_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08279__C _00896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07600_ _00216_ _04843_ _04907_ _00217_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a22o_1
XMuI._6474_ MuI._2340_ MuI._2362_ vssd1 vssd1 vccd1 vccd1 MuI._2365_ sky130_fd_sc_hd__and2_1
XANTENNA__13482__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3686_ MuI._2785_ vssd1 vssd1 vccd1 vccd1 MuI._2786_ sky130_fd_sc_hd__clkbuf_4
X_08580_ _01196_ _01197_ _01182_ _01184_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a211o_1
XFILLER_19_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5425_ MuI._1207_ MuI._1209_ MuI._1210_ vssd1 vssd1 vccd1 vccd1 MuI._1211_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07480__A _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07531_ _06659_ _06660_ _06673_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__nand3_1
XANTENNA__12098__A _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08295__B _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5356_ MuI._1132_ MuI._1133_ MuI._1134_ vssd1 vssd1 vccd1 vccd1 MuI._1135_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08726__D net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07462_ net118 net117 _04434_ _04509_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__and4_1
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11433__C _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4307_ MuI._3401_ MuI._3405_ vssd1 vssd1 vccd1 vccd1 MuI._3407_ sky130_fd_sc_hd__nand2_1
X_09201_ _06469_ _02194_ _04767_ net10 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__and4_1
XFILLER_167_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11208__B1 _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5287_ MuI._1057_ MuI._1058_ vssd1 vssd1 vccd1 vccd1 MuI._1059_ sky130_fd_sc_hd__or2b_1
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07393_ _06599_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__buf_6
XFILLER_176_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4238_ MuI._3332_ MuI._3336_ MuI._3325_ MuI._3337_ vssd1 vssd1 vccd1 vccd1 MuI._3338_
+ sky130_fd_sc_hd__o211ai_4
X_09132_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__or2_1
XANTENNA__11730__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06824__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4169_ MuI._3268_ vssd1 vssd1 vccd1 vccd1 MuI._3269_ sky130_fd_sc_hd__clkbuf_4
X_09063_ _01332_ _02334_ _00032_ _04767_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__and4_1
XFILLER_175_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07639__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08014_ _00623_ _00628_ _00624_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__nand3_1
XANTENNA__08461__D _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1406__D AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._766__B AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._485__C AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _02608_ _02624_ _02627_ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__o211ai_1
XANTENNA_MuI._4850__A2_N MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10081__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08916_ _01288_ _01285_ _01287_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__nand3_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09896_ _02302_ _03928_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__nand2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10498__A1 _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5303__B MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__B2 _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__nor2_1
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13436__A1 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07917__A2_N _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ _03002_ _00303_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__nand2_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13436__B2 _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0878__B_N net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__A _01096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _00281_ _03443_ _04240_ _04305_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__nand4_1
XANTENNA_MuI._6027__A1 MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6027__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10740_ _03460_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nand3_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ _03184_ _03188_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__nand2_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _02796_ _02792_ _02799_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21oi_1
XFILLER_167_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _02645_ _02694_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._3774__A MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _02984_ _06477_ _06546_ _03389_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__a22o_1
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6150__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10256__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12272_ _05109_ _05110_ _05092_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a21oi_2
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _03980_ _03981_ _03796_ _03799_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__o211a_1
XFILLER_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1650_ AuI._0606_ AuI._0004_ AuI._0005_ vssd1 vssd1 vccd1 vccd1 AuI.result\[25\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09764__B _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__A _05308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12902__C _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11154_ _02496_ _05895_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__nand2_1
XAuI._1581_ AuI._0633_ AuI._0754_ vssd1 vssd1 vccd1 vccd1 AuI._0756_ sky130_fd_sc_hd__and2b_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10105_ _03346_ _05467_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__and2b_1
X_11085_ _03691_ _03833_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__o21a_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10036_ net4 net3 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__or2b_1
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3540_ MuI.b_operand\[16\] vssd1 vssd1 vccd1 vccd1 MuI._1296_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._6028__C MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13427__A1 _02815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06909__A _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3471_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._0537_ sky130_fd_sc_hd__buf_2
XFILLER_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11438__B1 _04076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3949__A MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5210_ MuI._0883_ MuI._0884_ MuI._0894_ vssd1 vssd1 vccd1 vccd1 MuI._0974_ sky130_fd_sc_hd__a21oi_1
X_11987_ _04770_ _04804_ _04805_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__nor3_1
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6190_ MuI._2813_ MuI._2066_ MuI._2916_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._2052_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10938_ _02350_ _02742_ _02943_ _04133_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__a22o_1
XANTENNA__08854__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12650__A2 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5141_ MuI._2866_ MuI._2868_ MuI.a_operand\[8\] MuI.a_operand\[7\] vssd1 vssd1
+ vccd1 vccd1 MuI._0898_ sky130_fd_sc_hd__and4_1
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1015_ AuI._0199_ AuI._0200_ AuI._0226_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0227_
+ sky130_fd_sc_hd__a31oi_1
XFILLER_189_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ _06598_ _06599_ _06489_ _05498_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__and4_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5072_ MuI._2850_ MuI._0315_ MuI._0820_ MuI._0821_ vssd1 vssd1 vccd1 vccd1 MuI._0822_
+ sky130_fd_sc_hd__a31o_1
X_13037__134 vssd1 vssd1 vccd1 vccd1 _13037__134/HI net134 sky130_fd_sc_hd__conb_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _05471_ _05472_ _05329_ _05331_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__o211a_1
XANTENNA_MuI._5883__B MuI._1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12402__A2 _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__C net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4023_ MuI._3085_ MuI._3086_ MuI._3121_ MuI._3122_ vssd1 vssd1 vccd1 vccd1 MuI._3123_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11610__B1 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ _05154_ _05268_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__or2_1
XANTENNA__10166__A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10964__A2 _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5974_ MuI._1812_ MuI._1814_ vssd1 vssd1 vccd1 vccd1 MuI._1815_ sky130_fd_sc_hd__and2_1
XFILLER_125_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5107__C MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0969__A0 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4925_ MuI._0659_ MuI._0660_ vssd1 vssd1 vccd1 vccd1 MuI._0661_ sky130_fd_sc_hd__nor2_1
XANTENNA__12812__C _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07475__A _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11709__B _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._785_ AuI.pe._319_ AuI.pe._323_ AuI.pe._324_ AuI.pe._325_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._326_ sky130_fd_sc_hd__or4_1
XMuI._4856_ MuI._0572_ MuI._0573_ MuI._0584_ vssd1 vssd1 vccd1 vccd1 MuI._0585_ sky130_fd_sc_hd__nand3_2
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09750_ _02219_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__xnor2_1
X_06962_ net13 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__clkbuf_8
XFILLER_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3807_ MuI._2066_ MuI._2850_ vssd1 vssd1 vccd1 vccd1 MuI._2907_ sky130_fd_sc_hd__nand2_1
XFILLER_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08701_ _01202_ _01317_ _01318_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__and3_1
XMuI._4787_ MuI._0379_ MuI._0508_ vssd1 vssd1 vccd1 vccd1 MuI._0509_ sky130_fd_sc_hd__nor2_1
X_09681_ _02317_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__or2_1
X_06893_ _04273_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_55_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6526_ MuI._2420_ MuI._2415_ MuI._2419_ vssd1 vssd1 vccd1 vccd1 MuI._2422_ sky130_fd_sc_hd__and3_1
XMuI._3738_ MuI._2837_ vssd1 vssd1 vccd1 vccd1 MuI._2838_ sky130_fd_sc_hd__buf_2
X_08632_ _00444_ _00301_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4268__B1 MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06819__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6457_ MuI._1950_ MuI._1953_ MuI._1951_ vssd1 vssd1 vccd1 vccd1 MuI._2346_ sky130_fd_sc_hd__o21ba_1
XMuI._3669_ MuI._2627_ MuI._2649_ MuI._2682_ MuI._2704_ vssd1 vssd1 vccd1 vccd1 MuI._2715_
+ sky130_fd_sc_hd__a22o_1
X_08563_ _00934_ _00935_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__xor2_1
XFILLER_208_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09098__A1 _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09098__B2 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5408_ MuI._1134_ MuI._1132_ MuI._1133_ vssd1 vssd1 vccd1 vccd1 MuI._1192_ sky130_fd_sc_hd__or3_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ net117 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__buf_4
XMuI._6388_ MuI._2083_ MuI._2084_ MuI._2098_ vssd1 vssd1 vccd1 vccd1 MuI._2270_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08494_ _01108_ _01109_ _01111_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__o21a_1
XFILLER_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08845__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5339_ MuI._1108_ MuI._1113_ MuI._1114_ MuI._1115_ vssd1 vssd1 vccd1 vccd1 MuI._1116_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07445_ _00028_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__buf_4
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07376_ _06675_ _06674_ _06642_ _06556_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__o211a_1
XFILLER_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09115_ _01611_ _01613_ _01614_ _01381_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_148_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11092__A1_N _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10955__A2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _01644_ _01645_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__or4bb_1
XFILLER_191_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07385__A _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10523__B _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5314__A MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09948_ _02598_ _02600_ _02601_ _02602_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a211oi_1
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6248__A1 MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _02259_ _03982_ _02493_ _02494_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__o2bb2a_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _04533_ _04541_ _04540_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o21bai_1
XFILLER_46_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12890_ _02809_ _05773_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__nand2_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3769__A MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _02871_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__xor2_1
XFILLER_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1137__A0 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5471__A2 MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3482__A1 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _00289_ _05036_ _05112_ _00290_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22o_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10643__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ _02345_ _02377_ _03444_ _05948_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__and4_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__B1 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10643__B2 _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08663__B _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ _03165_ _03169_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a211o_1
X_13442_ _06276_ _06285_ _06324_ _06325_ _06326_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__a32o_1
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13373_ _06276_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nand2_1
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ _02703_ _03295_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__xnor2_2
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4734__A1 MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4734__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12255_ _04919_ _04922_ _04920_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__o21bai_1
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ _00077_ _00550_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__nand2_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1633_ AuI._0686_ AuI._0690_ vssd1 vssd1 vccd1 vccd1 AuI._0798_ sky130_fd_sc_hd__xor2_1
X_12186_ _02795_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__or2_1
XMuI._4710_ MuI._2803_ MuI._2352_ MuI._2374_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._0424_
+ sky130_fd_sc_hd__a22oi_1
XMuI._5690_ MuI._1480_ MuI._1481_ MuI._1500_ MuI._1501_ vssd1 vssd1 vccd1 vccd1 MuI._1502_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11137_ _03718_ _03720_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__nand2_1
XAuI._1564_ AuI._0667_ AuI._0741_ vssd1 vssd1 vccd1 vccd1 AuI._0742_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._570_ AuI.pe._125_ AuI.pe._026_ AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 AuI.pe._126_
+ sky130_fd_sc_hd__a21o_1
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6039__B MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4641_ MuI._0169_ MuI._0347_ vssd1 vssd1 vccd1 vccd1 MuI._0348_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11068_ _03639_ _03641_ _03814_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__o211a_1
XAuI._1495_ AuI._0679_ AuI._0680_ vssd1 vssd1 vccd1 vccd1 AuI._0681_ sky130_fd_sc_hd__nand2_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12880__A2_N _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__A1 _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4572_ MuI._0270_ MuI._0271_ vssd1 vssd1 vccd1 vccd1 MuI._0272_ sky130_fd_sc_hd__xor2_1
XFILLER_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10019_ _02685_ _02686_ _02635_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o21a_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12320__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6311_ MuI._2161_ MuI._2162_ MuI._2184_ vssd1 vssd1 vccd1 vccd1 MuI._2185_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3523_ MuI._1087_ MuI._1098_ vssd1 vssd1 vccd1 vccd1 MuI._1109_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6242_ MuI._2814_ MuI._2813_ MuI._1021_ MuI._1483_ vssd1 vssd1 vccd1 vccd1 MuI._2109_
+ sky130_fd_sc_hd__and4_1
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3454_ MuI._0339_ vssd1 vssd1 vccd1 vccd1 MuI._0350_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07180__D _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6173_ MuI._2023_ MuI._2031_ MuI._2032_ vssd1 vssd1 vccd1 vccd1 MuI._2034_ sky130_fd_sc_hd__nand3_1
XFILLER_177_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5124_ MuI._0876_ MuI._0877_ MuI._0872_ vssd1 vssd1 vccd1 vccd1 MuI._0880_ sky130_fd_sc_hd__a21o_1
X_07230_ _06524_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10608__B _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5055_ MuI._0802_ MuI._0803_ vssd1 vssd1 vccd1 vccd1 MuI._0804_ sky130_fd_sc_hd__nor2_1
XFILLER_201_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _06460_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__nand2_1
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07189__B _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4303__A MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4006_ MuI._1153_ MuI._2528_ MuI._2797_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._3106_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5118__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _06397_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5957_ MuI._1777_ MuI._1779_ MuI._0730_ vssd1 vssd1 vccd1 vccd1 MuI._1796_ sky130_fd_sc_hd__o21ai_1
XANTENNA_MuI._3861__B MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4908_ MuI._0640_ MuI._0641_ MuI._2817_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._0642_
+ sky130_fd_sc_hd__and4bb_1
X_09802_ _06504_ net132 net127 _06503_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22oi_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5888_ MuI._1581_ MuI._1668_ MuI._1679_ MuI._1680_ vssd1 vssd1 vccd1 vccd1 MuI._1720_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07994_ _00610_ _00611_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__and2_1
XFILLER_87_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._768_ AuI.pe._089_ AuI.pe._304_ AuI.pe._309_ AuI.pe._311_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._312_ sky130_fd_sc_hd__a211o_1
XMuI._4839_ MuI._0562_ MuI._0565_ vssd1 vssd1 vccd1 vccd1 MuI._0566_ sky130_fd_sc_hd__nor2_1
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ _02370_ _02371_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__and2_1
X_06945_ _04832_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08748__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1367__A0 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._699_ AuI.pe._380_ AuI.pe._391_ AuI.pe._118_ AuI.pe._105_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._246_ sky130_fd_sc_hd__a22o_1
XANTENNA__11455__A _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09664_ _02277_ _02281_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__xnor2_1
X_06876_ net126 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__buf_2
XANTENNA__07869__A2 _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._6509_ MuI._1912_ MuI._2110_ vssd1 vssd1 vccd1 vccd1 MuI._2403_ sky130_fd_sc_hd__and2_1
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10873__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ _06593_ _04649_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__nand2_2
X_09595_ _06520_ _06516_ _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__and4_1
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10873__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _01161_ _01163_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__and2b_1
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3739__D MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11822__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _00913_ _00912_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__and2b_1
XANTENNA__08294__A2 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ net44 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__buf_4
XFILLER_211_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__B _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ _06656_ _06658_ _06657_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4213__A MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__A _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ _00762_ _00764_ _03063_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a211oi_1
XFILLER_164_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09029_ _01255_ _01571_ _01572_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__or3_1
XFILLER_191_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4716__B2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12040_ _04860_ _04861_ _04766_ _04746_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__o211ai_2
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4586__C MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07265__D _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__C net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12942_ _05829_ _05830_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__or2_1
XAuI._1280_ AuI._0429_ AuI._0447_ AuI._0479_ vssd1 vssd1 vccd1 vccd1 AuI._0480_ sky130_fd_sc_hd__nand3b_1
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07281__C _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _02039_ _05755_ _03314_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21a_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _02669_ _02724_ _04626_ _04630_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__a211o_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _03539_ _00678_ _06603_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__and3_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12627__C _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _06682_ _03424_ _03425_ _00000_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a22o_1
XFILLER_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07493__B1 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11686_ _04480_ _04481_ _04361_ _04362_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o211a_1
XFILLER_202_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ _06337_ _06339_ _04635_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__mux2_1
XFILLER_186_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _03339_ _03340_ _03350_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4123__A MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13356_ _04161_ _06258_ _06259_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a31o_1
X_10568_ _03043_ _03103_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06922__A _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0995_ AuI._0143_ AuI._0146_ vssd1 vssd1 vccd1 vccd1 AuI._0207_ sky130_fd_sc_hd__nand2_2
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6860_ MuI.b_operand\[23\] MuI._2489_ vssd1 vssd1 vccd1 vccd1 MuI._2763_ sky130_fd_sc_hd__nand2_1
XANTENNA__13318__B1 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12307_ _03013_ _05831_ _05043_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__and3_1
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _00921_ _01206_ _04907_ _04972_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__nand4_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10444__A _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ _06134_ _06195_ _06164_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and3_1
XMuI._5811_ MuI._1545_ MuI._1547_ MuI._1633_ MuI._1634_ vssd1 vssd1 vccd1 vccd1 MuI._1635_
+ sky130_fd_sc_hd__a211o_1
XMuI._6791_ MuI._2577_ MuI._2580_ vssd1 vssd1 vccd1 vccd1 MuI._2713_ sky130_fd_sc_hd__xnor2_1
X_12238_ _04977_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__inv_2
XMuI._5742_ MuI._1274_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._1559_ sky130_fd_sc_hd__nand2_1
XAuI._1616_ AuI._0693_ AuI._0781_ AuI._0784_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0785_
+ sky130_fd_sc_hd__o22a_1
X_12169_ _04998_ _05000_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__a21oi_1
XAuI.pe._622_ AuI.pe._033_ AuI.pe._142_ AuI.pe._395_ vssd1 vssd1 vccd1 vccd1 AuI.pe._174_
+ sky130_fd_sc_hd__and3_1
XFILLER_123_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11567__A1_N _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5673_ MuI.b_operand\[11\] MuI._2829_ vssd1 vssd1 vccd1 vccd1 MuI._1484_ sky130_fd_sc_hd__nand2_1
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1547_ AuI._0650_ AuI._0727_ vssd1 vssd1 vccd1 vccd1 AuI._0728_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._553_ AuI.pe._056_ AuI.pe._066_ AuI.pe._054_ AuI.pe._063_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._110_ sky130_fd_sc_hd__a22o_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4624_ MuI._0327_ MuI._2854_ MuI._2484_ MuI._2853_ vssd1 vssd1 vccd1 vccd1 MuI._0330_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_AuI._1349__B1 AuI._0542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 a_operand[0] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06730_ net106 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__buf_6
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3694__A1 MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1478_ AuI._0638_ AuI._0639_ vssd1 vssd1 vccd1 vccd1 AuI._0664_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4891__B1 MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._484_ AuI.pe._046_ AuI.pe._038_ vssd1 vssd1 vccd1 vccd1 AuI.pe._047_ sky130_fd_sc_hd__nand2_1
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4555_ MuI._0226_ MuI._0253_ vssd1 vssd1 vccd1 vccd1 MuI._0254_ sky130_fd_sc_hd__or2_1
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3506_ MuI._0812_ MuI._0823_ MuI._0834_ vssd1 vssd1 vccd1 vccd1 MuI._0922_ sky130_fd_sc_hd__o21ba_1
XFILLER_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08400_ _01016_ _01015_ _01003_ _00986_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__o211a_1
XMuI._4486_ MuI._0176_ MuI._0177_ vssd1 vssd1 vccd1 vccd1 MuI._0178_ sky130_fd_sc_hd__and2_1
XANTENNA__12057__B1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _06579_ _04100_ _00271_ _06578_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22oi_1
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6225_ MuI._2087_ MuI._2090_ vssd1 vssd1 vccd1 vccd1 MuI._2091_ sky130_fd_sc_hd__nor2_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3437_ MuI.a_operand\[28\] MuI.b_operand\[28\] vssd1 vssd1 vccd1 vccd1 MuI._0163_
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08331_ _00946_ _00945_ _00944_ _00908_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__o211a_1
XFILLER_178_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09473__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6156_ MuI._0779_ MuI._2550_ MuI._2517_ MuI._2894_ vssd1 vssd1 vccd1 vccd1 MuI._2015_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _00875_ _00876_ _00879_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__a21bo_1
XFILLER_178_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5107_ MuI._2785_ MuI._2341_ MuI._2885_ MuI._3307_ vssd1 vssd1 vccd1 vccd1 MuI._0861_
+ sky130_fd_sc_hd__and4_1
XFILLER_119_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ _02420_ _06513_ _05176_ _05241_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__and4_1
XFILLER_193_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6087_ MuI._1927_ MuI._1928_ MuI._1938_ vssd1 vssd1 vccd1 vccd1 MuI._1939_ sky130_fd_sc_hd__a21o_1
X_08193_ _00525_ _00526_ _00524_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a21boi_4
XFILLER_193_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_A net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5038_ MuI._0285_ MuI._0417_ vssd1 vssd1 vccd1 vccd1 MuI._0785_ sky130_fd_sc_hd__nor2_1
XFILLER_119_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07144_ _06442_ _03960_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__a22o_1
XANTENNA__09776__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06832__A _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__C _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07075_ _06222_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10354__A _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11169__B _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__C _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11335__A2 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08200__A2 _00663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07663__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _00096_ _04294_ _04358_ _00095_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__a22oi_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10801__B _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ _06492_ _06463_ _00266_ _00592_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__nand4_1
X_06928_ _04649_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__buf_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11616__C _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _02169_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__or2_1
X_06859_ _03906_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__buf_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4208__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11913__A _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09578_ _02170_ _02185_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__B _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08529_ _03217_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08267__A2 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__A2 _02875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10074__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _02786_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__inv_2
XANTENNA__11271__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ _04184_ _04185_ _04248_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__a211o_2
XFILLER_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12744__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._095_ FuI._055_ vssd1 vssd1 vccd1 vccd1 FuI._056_ sky130_fd_sc_hd__clkbuf_2
X_10422_ _03118_ _03120_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__nor2_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__B1 _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ _03755_ _05713_ _06115_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__a21o_1
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09767__A2 _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06742__A _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3782__A MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10353_ _05305_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__buf_4
X_13141_ _06042_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__nor2_1
XFILLER_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07557__B _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _03809_ _05520_ _05969_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__nand3_1
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input56_A b_operand[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _02960_ _02961_ _02972_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12023_ _04831_ _04842_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__and3_1
XFILLER_133_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1401_ AuI._0581_ AuI._0573_ AuI._0590_ vssd1 vssd1 vccd1 vccd1 AuI._0591_ sky130_fd_sc_hd__a21o_1
XANTENNA__07573__A _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1332_ AuI._0526_ AuI._0527_ vssd1 vssd1 vccd1 vccd1 AuI._0528_ sky130_fd_sc_hd__xor2_2
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5221__B MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _05811_ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__nand2_1
XAuI._1263_ AuI._0448_ AuI._0451_ AuI._0463_ vssd1 vssd1 vccd1 vccd1 AuI._0464_ sky130_fd_sc_hd__a21o_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12919__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4340_ MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 MuI._0018_ sky130_fd_sc_hd__buf_2
XFILLER_73_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1194_ AuI._0328_ AuI._0326_ AuI._0347_ AuI._0348_ AuI._0399_ vssd1 vssd1 vccd1
+ vccd1 AuI._0400_ sky130_fd_sc_hd__o311ai_2
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ _05655_ _05658_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__A _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12638__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4271_ MuI.a_operand\[3\] vssd1 vssd1 vccd1 vccd1 MuI._3371_ sky130_fd_sc_hd__clkbuf_4
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _04480_ _04482_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__nor2_1
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08258__A2 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6010_ MuI._2550_ MuI._2517_ MuI._2066_ MuI._2916_ vssd1 vssd1 vccd1 vccd1 MuI._1854_
+ sky130_fd_sc_hd__and4_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _05559_ _05561_ _05663_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__a211oi_2
XFILLER_202_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__C _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11738_ _04534_ _04535_ _04536_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10158__B _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11669_ _04283_ _04447_ _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o211ai_2
X_13408_ _06320_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ _06191_ _06192_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nand2_1
XANTENNA__10174__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0978_ AuI._0154_ AuI._0162_ vssd1 vssd1 vccd1 vccd1 AuI._0190_ sky130_fd_sc_hd__xor2_2
XANTENNA__10773__B1 _03496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6843_ MuI._2753_ vssd1 vssd1 vccd1 vccd1 MuI.result\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6774_ MuI._2680_ MuI._2684_ MuI._2690_ MuI._2692_ MuI._2694_ vssd1 vssd1 vccd1
+ vccd1 MuI._2695_ sky130_fd_sc_hd__o2111a_1
XFILLER_102_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ _00503_ _00517_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__xnor2_4
XMuI._3986_ MuI._3011_ MuI._3025_ vssd1 vssd1 vccd1 vccd1 MuI._3086_ sky130_fd_sc_hd__or2b_1
X_08880_ _01449_ _01450_ _01451_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__o21ba_1
XMuI._5725_ MuI._1048_ MuI._1504_ MuI._1539_ MuI._1540_ vssd1 vssd1 vccd1 vccd1 MuI._1541_
+ sky130_fd_sc_hd__a211o_1
XFILLER_111_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07831_ _00221_ _04854_ _00446_ _00447_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__nand4_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11717__B _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._605_ AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 AuI.pe._158_ sky130_fd_sc_hd__buf_2
XANTENNA__07914__C _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08298__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5656_ MuI._1057_ MuI._1058_ MuI._0992_ vssd1 vssd1 vccd1 vccd1 MuI._1465_ sky130_fd_sc_hd__and3b_1
XFILLER_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ _00377_ _00378_ _00379_ vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__nand3_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._536_ AuI.pe._029_ AuI.pe._086_ AuI.pe._093_ vssd1 vssd1 vccd1 vccd1 AuI.pe._094_
+ sky130_fd_sc_hd__a21o_1
XMuI._4607_ MuI._0232_ MuI._0310_ vssd1 vssd1 vccd1 vccd1 MuI._0311_ sky130_fd_sc_hd__xnor2_1
X_09501_ _02124_ _02126_ _02125_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a21o_1
XMuI._5587_ MuI._1386_ MuI._1387_ MuI._1388_ vssd1 vssd1 vccd1 vccd1 MuI._1389_ sky130_fd_sc_hd__o21bai_1
XANTENNA_MuI._5131__B MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06713_ _02334_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__buf_4
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07693_ _00279_ _06436_ _04035_ _03378_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4028__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._467_ AuI.pe._029_ AuI.pe._020_ AuI.pe._031_ vssd1 vssd1 vccd1 vccd1 AuI.pe._032_
+ sky130_fd_sc_hd__o21a_1
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4538_ MuI._0099_ MuI._0234_ vssd1 vssd1 vccd1 vccd1 MuI._0235_ sky130_fd_sc_hd__xnor2_1
X_09432_ _02442_ _02496_ _00272_ _00301_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__and4_1
XFILLER_198_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06827__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._4970__B MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3867__A MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4588__A2_N MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4469_ MuI._0157_ MuI._0158_ vssd1 vssd1 vccd1 vccd1 MuI._0159_ sky130_fd_sc_hd__or2_1
X_09363_ _01965_ _01979_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__nand3_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4092__B2 MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6208_ MuI._2043_ MuI._2045_ MuI._2062_ vssd1 vssd1 vccd1 vccd1 MuI._2072_ sky130_fd_sc_hd__o21ai_1
XFILLER_178_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07457__B1 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _00915_ _00930_ _00931_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _01906_ _01910_ _01898_ _01911_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o211ai_1
XFILLER_20_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6139_ MuI._1994_ MuI._1995_ vssd1 vssd1 vccd1 vccd1 MuI._1996_ sky130_fd_sc_hd__nor2_1
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08245_ _00539_ _00836_ _00837_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__or3_1
XANTENNA__08761__B _01378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _00792_ _00793_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__xnor2_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07127_ _06427_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__clkbuf_8
XFILLER_133_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13098__C _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10084__A _01988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _06045_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4848__D MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11308__A2 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13395__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__B _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07393__A _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1441__B AuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4864__C MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07543__D net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10971_ _03708_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__xnor2_4
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _05581_ _02856_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__or2b_1
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11492__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11492__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06737__A _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _05416_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__or2_1
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5695__C MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10259__A _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3496__B MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _05423_ _05424_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07999__A1 _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12992__A1 _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__B2 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _04304_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__nand2_1
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._147_ FuI._009_ net153 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[18\] sky130_fd_sc_hd__dlxtn_1
XFILLER_184_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0901_ AuI._0119_ AuI._0120_ vssd1 vssd1 vccd1 vccd1 AuI._0121_ sky130_fd_sc_hd__nor2_1
X_11454_ _00878_ _05702_ _05767_ _00877_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__a22oi_1
XFILLER_172_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._078_ FuI._035_ FuI._043_ FuI.a_operand\[3\] vssd1 vssd1 vccd1 vccd1 FuI._015_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11547__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0832_ AuI._0050_ net124 net125 AuI._0051_ vssd1 vssd1 vccd1 vccd1 AuI._0052_
+ sky130_fd_sc_hd__a22o_1
X_10405_ _03100_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__xor2_2
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11385_ _02709_ _02064_ _06023_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or3b_1
XFILLER_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _06024_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__nand2_1
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10336_ _03163_ _04789_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__and2_1
XANTENNA__07620__B1 _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3840_ MuI._1142_ MuI._2495_ MuI._2791_ MuI._2939_ vssd1 vssd1 vccd1 vccd1 MuI._2940_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11818__A _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _00672_ _00711_ _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__o21ai_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _05867_ _05874_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a21o_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10722__A _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3771_ MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 MuI._2871_ sky130_fd_sc_hd__clkbuf_4
X_12006_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__and2_1
XFILLER_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _04133_ _02302_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__or2b_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5510_ MuI._1255_ MuI._1254_ MuI._1253_ vssd1 vssd1 vccd1 vccd1 MuI._1304_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6490_ MuI._1917_ MuI._1992_ MuI._1990_ vssd1 vssd1 vccd1 vccd1 MuI._2382_ sky130_fd_sc_hd__a21oi_2
XFILLER_78_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5441_ MuI._1156_ MuI._1165_ MuI._1163_ vssd1 vssd1 vccd1 vccd1 MuI._1228_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._6047__B MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1315_ AuI._0509_ AuI._0512_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[14\]
+ sky130_fd_sc_hd__xnor2_4
XFILLER_207_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08846__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5372_ MuI._1139_ MuI._1150_ MuI._1151_ vssd1 vssd1 vccd1 vccd1 MuI._1152_ sky130_fd_sc_hd__nand3_1
XFILLER_207_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ _05793_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__and2_1
XFILLER_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1246_ AuI._0344_ AuI._0413_ AuI._0442_ vssd1 vssd1 vccd1 vccd1 AuI._0448_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._5886__B MuI._1662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4323_ MuI._3390_ MuI._3421_ MuI._3422_ vssd1 vssd1 vccd1 vccd1 MuI._0000_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3687__A MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11272__B _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__A1 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12839_ _05631_ _05634_ _05632_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__o21ba_1
XAuI._1177_ AuI._0177_ AuI._0188_ AuI._0311_ AuI._0183_ AuI._0208_ AuI._0307_ vssd1
+ vssd1 vccd1 vccd1 AuI._0383_ sky130_fd_sc_hd__mux4_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6063__A MuI._3154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__B2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4254_ MuI._3345_ MuI._3347_ vssd1 vssd1 vccd1 vccd1 MuI._3354_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08100__A1 _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4185_ MuI._3282_ MuI._3284_ vssd1 vssd1 vccd1 vccd1 MuI._3285_ sky130_fd_sc_hd__and2b_1
XANTENNA__10319__D _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4014__C MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08030_ _00579_ _00584_ _00564_ _00585_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__a211o_1
XANTENNA__07478__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 a_operand[3] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_4
Xinput41 b_operand[13] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_6
Xinput52 b_operand[23] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_4
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 b_operand[4] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_6
XFILLER_190_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08403__A2 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10335__C _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10210__A2 _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _01631_ _01852_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o211ai_2
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6826_ MuI._2702_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2745_ sky130_fd_sc_hd__and2b_1
X_08932_ _01521_ _01526_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__and2_1
XFILLER_170_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3969_ MuI._3067_ MuI._3068_ vssd1 vssd1 vccd1 vccd1 MuI._3069_ sky130_fd_sc_hd__nor2_1
XMuI._6757_ MuI._2643_ MuI._2647_ MuI._2675_ vssd1 vssd1 vccd1 vccd1 MuI._2676_ sky130_fd_sc_hd__nand3_1
X_08863_ _01470_ _01471_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__nand3_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10351__B _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__B1 _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5708_ MuI._1520_ MuI._1521_ vssd1 vssd1 vccd1 vccd1 MuI._1522_ sky130_fd_sc_hd__nor2_1
XFILLER_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6688_ MuI._2593_ MuI._2599_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2600_ sky130_fd_sc_hd__mux2_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07814_ _00428_ _00429_ _00410_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a21o_1
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08794_ _01410_ _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__or2_1
XFILLER_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5639_ MuI._1429_ MuI._1409_ MuI._1401_ vssd1 vssd1 vccd1 vccd1 MuI._1446_ sky130_fd_sc_hd__and3b_1
XANTENNA_MuI._4301__A2 MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07745_ _06458_ _00362_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__or2_1
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._519_ AuI.pe._078_ vssd1 vssd1 vccd1 vccd1 AuI.pe._079_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13463__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__B _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07676_ _00283_ _04046_ _00288_ _00291_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3597__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _01957_ _01924_ _01956_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__or3_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__A _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13215__A2 _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _01882_ _01883_ _01958_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a21o_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08772__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _01779_ _01888_ _01884_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__and3_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1494__A2 AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _00835_ _00844_ _00845_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__nand3_2
XFILLER_154_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08159_ _00775_ _00774_ _00773_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _03924_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _02916_ _04929_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__or2b_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10542__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _02722_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6148__A MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5052__A MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4828__B1 MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input19_A a_operand[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1100_ AuI._0269_ AuI._0267_ AuI._0176_ vssd1 vssd1 vccd1 vccd1 AuI._0310_ sky130_fd_sc_hd__mux2_1
XFILLER_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10954_ _03511_ _03655_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__nand2_1
XFILLER_204_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1031_ net110 net30 net59 net27 AuI._0123_ AuI._0174_ vssd1 vssd1 vccd1 vccd1
+ AuI._0243_ sky130_fd_sc_hd__mux4_1
XFILLER_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10885_ _03598_ _03617_ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__nand3_2
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12624_ _02856_ _05488_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
XANTENNA__09778__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12965__B2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12555_ _05039_ _05151_ _05415_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__o21ai_1
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4359__A2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11506_ _04285_ _04286_ _04127_ _04270_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a211o_1
XANTENNA__07298__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07729__C _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ _03842_ _04994_ _05216_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a31o_1
XFILLER_172_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12717__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5990_ MuI._1817_ MuI._1825_ MuI._1828_ MuI._1827_ vssd1 vssd1 vccd1 vccd1 MuI._1832_
+ sky130_fd_sc_hd__a211o_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _04076_ _04207_ _04212_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o211a_1
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4941_ MuI._0675_ MuI._0677_ vssd1 vssd1 vccd1 vccd1 MuI._0678_ sky130_fd_sc_hd__nor2_1
XANTENNA__12193__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__B1 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output87_A net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._0815_ AuI._0025_ net114 AuI._0028_ AuI._0033_ AuI._0034_ vssd1 vssd1 vccd1 vccd1
+ AuI._0035_ sky130_fd_sc_hd__o221a_1
XANTENNA__06930__A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11368_ _04094_ _04095_ _04138_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__and4_1
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4872_ MuI._0599_ MuI._0601_ vssd1 vssd1 vccd1 vccd1 MuI._0602_ sky130_fd_sc_hd__and2_1
X_13107_ _03489_ _06002_ _06005_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a211o_1
X_10319_ _02905_ _02959_ _00421_ _00423_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__nand4_1
XFILLER_140_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11299_ _04063_ _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__nand3_1
XMuI._3823_ MuI._2913_ MuI._2922_ vssd1 vssd1 vccd1 vccd1 MuI._2923_ sky130_fd_sc_hd__xor2_2
XMuI._6611_ MuI._1462_ MuI._1555_ MuI._1642_ vssd1 vssd1 vccd1 vccd1 MuI._2515_ sky130_fd_sc_hd__nor3b_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _03293_ _02724_ _05931_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__a211o_1
XANTENNA__11267__B _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10171__B _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6542_ MuI._2428_ MuI._2228_ vssd1 vssd1 vccd1 vccd1 MuI._2439_ sky130_fd_sc_hd__and2b_1
XFILLER_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3754_ MuI.b_operand\[9\] vssd1 vssd1 vccd1 vccd1 MuI._2854_ sky130_fd_sc_hd__buf_2
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08857__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6473_ MuI._2340_ MuI._2362_ vssd1 vssd1 vccd1 vccd1 MuI._2364_ sky130_fd_sc_hd__nor2_1
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3685_ MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 MuI._2785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5424_ MuI._2873_ MuI._2875_ MuI._0444_ MuI.a_operand\[1\] vssd1 vssd1 vccd1
+ vccd1 MuI._1210_ sky130_fd_sc_hd__and4_1
XFILLER_208_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07530_ _00026_ _00027_ _00146_ _00147_ vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__nand4_1
XFILLER_35_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12098__B _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5355_ MuI.a_operand\[8\] MuI.a_operand\[7\] MuI._3402_ MuI._3396_ vssd1 vssd1
+ vccd1 vccd1 MuI._1134_ sky130_fd_sc_hd__and4_1
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08295__C _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07461_ _00076_ _00078_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__nor2_1
XAuI._1229_ AuI._0429_ AuI._0432_ vssd1 vssd1 vccd1 vccd1 AuI._0433_ sky130_fd_sc_hd__and2_1
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4306_ MuI._3401_ MuI._3405_ vssd1 vssd1 vccd1 vccd1 MuI._3406_ sky130_fd_sc_hd__xor2_2
XANTENNA__11433__D _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ _06463_ _04767_ _06602_ _02107_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22oi_2
XMuI._5286_ MuI._1055_ MuI._1056_ MuI._0928_ MuI._0952_ vssd1 vssd1 vccd1 vccd1 MuI._1058_
+ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._6224__C MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11208__A1 _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07392_ _06606_ _06601_ _06584_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and3_1
XFILLER_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11208__B2 _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08232__A2_N _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4237_ MuI._3315_ MuI._3322_ MuI._3324_ vssd1 vssd1 vccd1 vccd1 MuI._3337_ sky130_fd_sc_hd__nand3_1
XFILLER_176_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09131_ _01737_ _01746_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__xor2_1
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__B _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4168_ MuI.b_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._3268_ sky130_fd_sc_hd__clkbuf_4
X_09062_ _01601_ _01598_ _01600_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__nand3_1
XANTENNA__10185__A_N _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07639__C _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08013_ _00529_ _00630_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07001__A _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4099_ MuI._2605_ MuI._2844_ MuI._2845_ MuI._2840_ vssd1 vssd1 vccd1 vccd1 MuI._3199_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_163_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__B1 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09964_ _02596_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__or2_1
XANTENNA_AuI.pe._485__D AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6809_ MuI._0086_ MuI._2732_ vssd1 vssd1 vccd1 vccd1 MuI._2733_ sky130_fd_sc_hd__xor2_4
XANTENNA__13133__A1 _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4522__A2 MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _01495_ _01496_ _01505_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__nand3_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09895_ _02543_ _02538_ _02542_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nor3_1
XANTENNA__10081__B _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08846_ _01332_ _02334_ _06602_ _06604_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__and4_1
XANTENNA__10498__A2 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07671__A _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08777_ _01359_ _01361_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__nor2_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13436__A2 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12289__A _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _03443_ _04240_ _04305_ _00290_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a22o_1
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6027__A2 MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11998__A2 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07659_ _00275_ _00276_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._4216__A MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10670_ _03384_ _03385_ _03381_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a21o_1
XFILLER_167_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _01898_ _01911_ _01906_ _01910_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a211o_1
XANTENNA__08076__B1 _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ _03335_ _05456_ _05055_ _05054_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a31o_1
XFILLER_166_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08007__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6150__B MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10256__B _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ _05092_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__and3_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._800__B1 AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11222_ _03796_ _03799_ _03980_ _03981_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a211oi_4
XANTENNA__07846__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1580_ AuI._0754_ AuI._0633_ vssd1 vssd1 vccd1 vccd1 AuI._0755_ sky130_fd_sc_hd__and2b_1
X_11153_ _03808_ _03799_ _03800_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__nand3_1
XANTENNA__12902__D _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _02777_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__nor2_1
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11084_ _03691_ _03833_ _06428_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10035_ net2 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11686__A1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08551__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6028__D MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3470_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._0526_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._3949__B MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__B1 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _04803_ _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__and3_1
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _02718_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08854__A2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5140_ MuI._0168_ MuI._2319_ vssd1 vssd1 vccd1 vccd1 MuI._0897_ sky130_fd_sc_hd__nand2_1
XANTENNA__12927__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1014_ net38 net6 AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0226_ sky130_fd_sc_hd__mux2_1
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _06630_ _05445_ _05509_ _06631_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__a22oi_1
XMuI._5071_ MuI._2853_ MuI._2854_ MuI.a_operand\[3\] MuI._0444_ vssd1 vssd1 vccd1
+ vccd1 MuI._0821_ sky130_fd_sc_hd__and4_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__A _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _05329_ _05331_ _05471_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a211oi_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4022_ MuI._3119_ MuI._3120_ MuI._3088_ MuI._3089_ vssd1 vssd1 vccd1 vccd1 MuI._3122_
+ sky130_fd_sc_hd__a211oi_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _03525_ _04316_ _03343_ _03342_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__a31o_1
XFILLER_158_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09658__D _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11610__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ _05222_ _05224_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__o211ai_4
XFILLER_172_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11610__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _05196_ _05199_ _05322_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o211ai_1
XANTENNA__12662__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07756__A _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5973_ MuI._1811_ MuI._1795_ MuI._1810_ vssd1 vssd1 vccd1 vccd1 MuI._1814_ sky130_fd_sc_hd__nand3_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5107__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4924_ MuI._0649_ MuI._0651_ MuI._0657_ vssd1 vssd1 vccd1 vccd1 MuI._0660_ sky130_fd_sc_hd__and3_1
XFILLER_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0969__A1 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12812__D _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._784_ AuI.pe._397_ AuI.pe._173_ vssd1 vssd1 vccd1 vccd1 AuI.pe._325_ sky130_fd_sc_hd__or2_1
XANTENNA_AuI._0827__A_N net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4855_ MuI._0577_ MuI._0583_ vssd1 vssd1 vccd1 vccd1 MuI._0584_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06961_ _05005_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[16\] sky130_fd_sc_hd__clkbuf_2
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3806_ MuI._2879_ MuI._2904_ MuI._2905_ vssd1 vssd1 vccd1 vccd1 MuI._2906_ sky130_fd_sc_hd__a21boi_2
X_08700_ _01188_ _01191_ _01190_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__o21ai_1
XMuI._4786_ MuI._1461_ MuI._0378_ MuI._0376_ MuI._0377_ vssd1 vssd1 vccd1 vccd1 MuI._0508_
+ sky130_fd_sc_hd__o2bb2a_1
X_09680_ _02319_ _02321_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__xnor2_2
XANTENNA_AuI.pe._570__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06892_ _04262_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__and3_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3737_ MuI.b_operand\[9\] vssd1 vssd1 vccd1 vccd1 MuI._2837_ sky130_fd_sc_hd__buf_2
XMuI._6525_ MuI._2415_ MuI._2419_ MuI._2420_ vssd1 vssd1 vccd1 vccd1 MuI._2421_ sky130_fd_sc_hd__a21o_1
XANTENNA__07491__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08631_ _01246_ _01248_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nor2_1
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3668_ MuI._2693_ vssd1 vssd1 vccd1 vccd1 MuI._2704_ sky130_fd_sc_hd__buf_2
XMuI._6456_ MuI._1949_ MuI._1954_ MuI._2344_ vssd1 vssd1 vccd1 vccd1 MuI._2345_ sky130_fd_sc_hd__a21oi_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ _01175_ _01178_ _01177_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__o21a_1
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09098__A2 _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5407_ MuI._1189_ MuI._1190_ vssd1 vssd1 vccd1 vccd1 MuI._1191_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6387_ MuI._2065_ MuI._2268_ vssd1 vssd1 vccd1 vccd1 MuI._2269_ sky130_fd_sc_hd__xor2_2
X_07513_ _00088_ _04520_ vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__nand2_1
XMuI._3599_ MuI._1923_ MuI._1934_ vssd1 vssd1 vccd1 vccd1 MuI._1945_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4036__A MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ _00918_ _01110_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08845__A2 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12837__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5338_ MuI._0978_ MuI._0980_ vssd1 vssd1 vccd1 vccd1 MuI._1115_ sky130_fd_sc_hd__and2_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07444_ _00029_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__buf_6
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06835__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3875__A MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5269_ MuI.a_operand\[15\] MuI.a_operand\[14\] MuI._0017_ MuI._0018_ vssd1 vssd1
+ vccd1 vccd1 MuI._1039_ sky130_fd_sc_hd__and4_1
XFILLER_22_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07375_ _06556_ _06642_ _06674_ _06675_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a211oi_4
XANTENNA__10357__A _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ _01711_ _01729_ _01730_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nor4_4
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3594__B MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09045_ _01644_ _01645_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13354__A1 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07385__B _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5314__B MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ _02601_ _02602_ _02598_ _02600_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__o211ai_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _02259_ _03895_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__and3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6248__A2 MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08829_ _01441_ _01445_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__nand3_1
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09105__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _02861_ _04624_ _01349_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__o21a_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12617__B1 _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1137__A1 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _04400_ _04404_ _04401_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__o21bai_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3482__A2 MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11651__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10722_ _00153_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__clkbuf_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10643__A2 _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06745__A _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09121__A _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ _02812_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _03366_ _03367_ _03356_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._6161__A MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _06283_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__inv_2
XFILLER_182_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08960__A _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10584_ _00814_ _03122_ _03123_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__o21a_1
XFILLER_139_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _03163_ _03449_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nand2_1
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4734__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12254_ _04923_ _04932_ _04931_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._3942__B1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11205_ _03962_ _03963_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._5505__A MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1632_ AuI._0259_ AuI._0796_ AuI._0797_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[20\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA_AuI._1073__A0 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ _05017_ _02897_ _02928_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1563_ AuI._0636_ AuI._0736_ vssd1 vssd1 vccd1 vccd1 AuI._0741_ sky130_fd_sc_hd__nor2_1
X_11136_ _03886_ _03887_ _03882_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a21o_1
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3670__D MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4640_ MuI._0171_ MuI._0170_ vssd1 vssd1 vccd1 vccd1 MuI._0347_ sky130_fd_sc_hd__nor2_1
XAuI._1494_ AuI._0375_ AuI._0498_ AuI._0577_ vssd1 vssd1 vccd1 vccd1 AuI._0680_ sky130_fd_sc_hd__o21bai_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11067_ _03776_ _03778_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__or4bb_2
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4571_ MuI._0112_ MuI._0471_ MuI._0109_ MuI._0107_ vssd1 vssd1 vccd1 vccd1 MuI._0271_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12320__A2 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _02635_ _02685_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__nor3_1
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._6310_ MuI._2169_ MuI._2183_ vssd1 vssd1 vccd1 vccd1 MuI._2184_ sky130_fd_sc_hd__xor2_1
XMuI._3522_ MuI._1043_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._1098_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4782__C MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6241_ MuI._2860_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._2108_ sky130_fd_sc_hd__nand2_1
XMuI._3453_ MuI._0328_ vssd1 vssd1 vccd1 vccd1 MuI._0339_ sky130_fd_sc_hd__clkbuf_4
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11969_ _03282_ _05380_ _05445_ _00124_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22oi_2
XANTENNA__12657__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6172_ MuI._2019_ MuI._2021_ MuI._2020_ vssd1 vssd1 vccd1 vccd1 MuI._2032_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13252__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5123_ MuI._0872_ MuI._0876_ MuI._0877_ vssd1 vssd1 vccd1 vccd1 MuI._0879_ sky130_fd_sc_hd__nand3_1
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5054_ MuI._2875_ MuI._3362_ MuI._0100_ MuI._2873_ vssd1 vssd1 vccd1 vccd1 MuI._0803_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07160_ net22 vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4005_ MuI._2814_ MuI._1142_ MuI._2528_ MuI._2539_ vssd1 vssd1 vccd1 vccd1 MuI._3105_
+ sky130_fd_sc_hd__and4_1
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _04929_ _06284_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__and2_1
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11347__B1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4957__C MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5956_ MuI._1768_ MuI._1794_ vssd1 vssd1 vccd1 vccd1 MuI._1795_ sky130_fd_sc_hd__nand2_1
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4907_ MuI._1153_ MuI._0111_ MuI._0315_ MuI._0735_ vssd1 vssd1 vccd1 vccd1 MuI._0641_
+ sky130_fd_sc_hd__a22oi_1
X_09801_ _02422_ _02421_ _02413_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a21o_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5887_ MuI._1164_ MuI._0421_ MuI._1663_ vssd1 vssd1 vccd1 vccd1 MuI._1719_ sky130_fd_sc_hd__and3_1
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07993_ _00600_ _00601_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__xnor2_1
XAuI.pe._767_ AuI.pe._380_ AuI.pe._395_ AuI.pe._310_ AuI.pe._132_ AuI.pe._378_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._311_ sky130_fd_sc_hd__a32o_1
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4838_ MuI._0563_ MuI._0564_ vssd1 vssd1 vccd1 vccd1 MuI._0565_ sky130_fd_sc_hd__or2_1
X_09732_ _02367_ _02369_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and2_1
XANTENNA__11736__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06944_ net10 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__buf_4
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._1367__A1 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._698_ AuI.pe._045_ AuI.pe._089_ AuI.pe._197_ AuI.pe._133_ AuI.pe._102_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._245_ sky130_fd_sc_hd__a32o_1
XANTENNA__08748__C _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4769_ MuI._0486_ MuI._0488_ vssd1 vssd1 vccd1 vccd1 MuI._0489_ sky130_fd_sc_hd__and2_1
X_09663_ _02289_ _02290_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__nand3_2
XANTENNA__11455__B _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _04079_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[2\] sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08110__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6508_ MuI._2213_ MuI._2226_ vssd1 vssd1 vccd1 vccd1 MuI._2402_ sky130_fd_sc_hd__nor2_1
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08614_ _01229_ _01231_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__nor2_1
X_09594_ _02229_ _04035_ _06433_ _02431_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22oi_2
XANTENNA__10873__A2 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6439_ MuI._2324_ MuI._2325_ vssd1 vssd1 vccd1 vccd1 MuI._2326_ sky130_fd_sc_hd__xnor2_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08545_ _01101_ _01162_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__nor2_1
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _03335_ _03982_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__nand2_1
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__B2 _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08483__C _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ _00028_ _00029_ _00035_ _04638_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__and4_1
XFILLER_211_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__C _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _06656_ _06657_ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nand3_2
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4213__B MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__B1 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__B _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07289_ _06583_ _05025_ _05112_ _06585_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__a22oi_1
XFILLER_191_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4716__A2 MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _01576_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__inv_2
XFILLER_164_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1444__B AuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4586__D MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11646__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__B _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10550__A _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _03831_ _05338_ _05728_ _05726_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a31oi_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _02039_ _05755_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__nand2_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07281__D _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11823_ FuI.Integer\[10\] _04627_ _03675_ _04671_ _04629_ vssd1 vssd1 vccd1 vccd1
+ _04630_ sky130_fd_sc_hd__a221o_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4942__A1_N MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11754_ _04464_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__inv_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10705_ _05627_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__clkbuf_4
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12627__D _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__A1 _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07493__B2 _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ _04361_ _04362_ _04480_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a211oi_1
XFILLER_81_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ _06338_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__clkinv_2
XFILLER_186_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10636_ _03339_ _03340_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13355_ _03314_ _06261_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI._1294__A0 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10567_ _03100_ _03102_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nor2_1
XFILLER_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0994_ AuI._0205_ vssd1 vssd1 vccd1 vccd1 AuI._0206_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13318__A1 _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _05046_ _05045_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__and2b_1
XANTENNA__13318__B2 _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _06134_ _06164_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__a21o_1
X_10498_ _01206_ _04907_ _04972_ _00921_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__a22o_1
XANTENNA__10444__B _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5810_ MuI._1631_ MuI._1632_ MuI._1573_ vssd1 vssd1 vccd1 vccd1 MuI._1634_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6790_ MuI._2568_ MuI._2571_ vssd1 vssd1 vccd1 vccd1 MuI._2712_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12237_ _05038_ _05074_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__xor2_1
XFILLER_123_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5741_ MuI._1495_ MuI._1496_ MuI._1492_ vssd1 vssd1 vccd1 vccd1 MuI._1558_ sky130_fd_sc_hd__o21bai_2
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1615_ AuI._0677_ AuI._0619_ vssd1 vssd1 vccd1 vccd1 AuI._0784_ sky130_fd_sc_hd__xor2_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12168_ _04998_ _05000_ _03134_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__o21ai_1
XAuI.pe._621_ AuI.pe._172_ vssd1 vssd1 vccd1 vccd1 AuI.pe._173_ sky130_fd_sc_hd__buf_2
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10552__A1 _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5672_ MuI._1025_ MuI._1026_ MuI._1024_ vssd1 vssd1 vccd1 vccd1 MuI._1482_ sky130_fd_sc_hd__a21bo_1
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _03525_ _04456_ _03699_ _03698_ _04596_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a32o_2
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1546_ AuI._0649_ AuI._0723_ AuI._0646_ vssd1 vssd1 vccd1 vccd1 AuI._0727_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10460__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ _01206_ _03425_ _05702_ _00921_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a22o_1
XAuI.pe._552_ AuI.pe._107_ AuI.pe._108_ vssd1 vssd1 vccd1 vccd1 AuI.pe._109_ sky130_fd_sc_hd__and2b_1
XMuI._4623_ MuI.b_operand\[10\] MuI._0327_ MuI._2837_ MuI.a_operand\[11\] vssd1 vssd1
+ vccd1 vccd1 MuI._0329_ sky130_fd_sc_hd__and4_1
XFILLER_77_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 a_operand[10] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_6
XFILLER_77_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6066__A MuI._1848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1477_ AuI._0652_ AuI._0657_ AuI._0660_ AuI._0661_ AuI._0662_ vssd1 vssd1 vccd1
+ vccd1 AuI._0663_ sky130_fd_sc_hd__a32oi_4
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11091__A1_N _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4554_ MuI._0226_ MuI._0227_ MuI._0252_ vssd1 vssd1 vccd1 vccd1 MuI._0253_ sky130_fd_sc_hd__nor3_1
XAuI.pe._483_ AuI.pe._045_ vssd1 vssd1 vccd1 vccd1 AuI.pe._046_ sky130_fd_sc_hd__buf_2
XANTENNA__09170__A1 _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3505_ MuI._0900_ vssd1 vssd1 vccd1 vccd1 MuI._0911_ sky130_fd_sc_hd__inv_2
XANTENNA__07181__B1 _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4485_ MuI._0158_ MuI._0160_ MuI._0175_ vssd1 vssd1 vccd1 vccd1 MuI._0177_ sky130_fd_sc_hd__or3_1
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12387__A _05232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6224_ MuI._2087_ MuI._2089_ MuI.b_operand\[20\] MuI._2682_ vssd1 vssd1 vccd1
+ vccd1 MuI._2090_ sky130_fd_sc_hd__and4bb_1
XMuI._3436_ MuI.a_operand\[29\] MuI.b_operand\[29\] vssd1 vssd1 vccd1 vccd1 MuI._0152_
+ sky130_fd_sc_hd__or2_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ _00939_ _00941_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__and2b_1
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09473__A2 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6155_ MuI._0559_ MuI._0768_ MuI._3000_ MuI._2754_ vssd1 vssd1 vccd1 vccd1 MuI._2014_
+ sky130_fd_sc_hd__and4_1
XFILLER_178_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08261_ _00877_ _00878_ _04649_ _04714_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__nand4_2
XMuI._5106_ MuI._3349_ MuI._2885_ MuI._3185_ MuI._3223_ vssd1 vssd1 vccd1 vccd1 MuI._0860_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_193_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6086_ MuI._1929_ MuI._1937_ vssd1 vssd1 vccd1 vccd1 MuI._1938_ sky130_fd_sc_hd__xnor2_1
X_07212_ net66 vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__buf_4
XFILLER_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4946__A2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ _00669_ _00809_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__xor2_4
XFILLER_193_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5037_ MuI._0672_ MuI._0782_ MuI._0783_ vssd1 vssd1 vccd1 vccd1 MuI._0784_ sky130_fd_sc_hd__o21a_1
XFILLER_195_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07143_ net112 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__buf_2
XANTENNA__07928__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout119_A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _04391_ _06067_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__and2_1
XANTENNA__08750__D _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10354__B _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07366__D _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5939_ MuI._0725_ MuI._0726_ MuI._0732_ vssd1 vssd1 vccd1 vccd1 MuI._1776_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._819_ AuI.pe._344_ AuI.pe._357_ vssd1 vssd1 vccd1 vccd1 AuI.pe._358_ sky130_fd_sc_hd__and2b_1
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07976_ _03152_ _00267_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__nand2_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ _00150_ net124 net123 _06469_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
XANTENNA__12296__A1 _02584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06927_ _04638_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__buf_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11616__D _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ _02669_ _03906_ _03993_ _02604_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22oi_1
XFILLER_83_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06858_ _03895_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__buf_4
XFILLER_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08775__A _01391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4208__B MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__B _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09577_ _02204_ _02208_ _02209_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a211oi_2
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _03152_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08528_ _03271_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__buf_4
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._1439__B AuI._0519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__A2 _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _01070_ _01075_ _01076_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__nand3_1
XFILLER_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _04247_ _04222_ _04223_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__and3_2
XFILLER_184_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12744__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._094_ FuI._036_ FuI._054_ vssd1 vssd1 vccd1 vccd1 FuI._055_ sky130_fd_sc_hd__nor2_1
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A1 _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _00666_ _00812_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07227__B2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _05950_ _05952_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and2_1
X_10352_ _02808_ _05262_ _05327_ _02765_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a22oi_4
XFILLER_192_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1028__A0 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _05966_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10283_ _02969_ _02971_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__xor2_1
XFILLER_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08727__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _04841_ _04839_ _04840_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nand3_2
XANTENNA_input49_A b_operand[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1400_ AuI._0567_ AuI._0578_ vssd1 vssd1 vccd1 vccd1 AuI._0590_ sky130_fd_sc_hd__or2b_1
XANTENNA__07573__B _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._507__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1331_ net12 net44 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0527_ sky130_fd_sc_hd__mux2_2
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12287__A1 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12924_ _03744_ _05456_ _05810_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a21o_1
XAuI._1262_ AuI._0462_ vssd1 vssd1 vccd1 vccd1 AuI._0463_ sky130_fd_sc_hd__inv_2
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07933__A1_N _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__B1 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4118__B MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12919__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13236__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1193_ AuI._0362_ AuI._0363_ AuI._0379_ AuI._0380_ vssd1 vssd1 vccd1 vccd1 AuI._0399_
+ sky130_fd_sc_hd__and4b_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12855_ _05737_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__and2_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4270_ MuI._3368_ MuI._3369_ vssd1 vssd1 vccd1 vccd1 MuI._3370_ sky130_fd_sc_hd__nor2_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._150__156 vssd1 vssd1 vccd1 vccd1 FuI._150__156/HI net156 sky130_fd_sc_hd__conb_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _04610_ _04611_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__nand2_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12000__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _05663_ _05664_ _05559_ _05561_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__o211a_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11737_ _04534_ _04535_ _04536_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__or3_1
XANTENNA__12357__D _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A2 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _04460_ _04461_ _04278_ _04282_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06933__A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _03680_ _05992_ _02820_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__and3_1
X_10619_ _03820_ _04133_ _03155_ _03153_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a31o_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10455__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _00063_ _00216_ _05574_ _03425_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__nand4_1
XFILLER_128_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13338_ _06248_ _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__xor2_1
XFILLER_115_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10174__B _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0977_ AuI._0031_ vssd1 vssd1 vccd1 vccd1 AuI._0189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_143_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6842_ MuI._2723_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2753_ sky130_fd_sc_hd__and2b_1
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ _06176_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nand2_1
XFILLER_170_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6773_ MuI._2632_ MuI._2636_ vssd1 vssd1 vccd1 vccd1 MuI._2694_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07764__A _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3985_ MuI._3008_ MuI._3010_ vssd1 vssd1 vccd1 vccd1 MuI._3085_ sky130_fd_sc_hd__or2_1
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5724_ MuI._1536_ MuI._1537_ MuI._1518_ vssd1 vssd1 vccd1 vccd1 MuI._1540_ sky130_fd_sc_hd__a21oi_1
X_07830_ _00444_ _00445_ _00446_ _00447_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a22o_1
XFILLER_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._604_ AuI.pe._102_ AuI.pe._066_ AuI.pe._054_ AuI.pe._106_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._157_ sky130_fd_sc_hd__a22o_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11717__C _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07914__D _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5655_ MuI._0844_ MuI._1061_ MuI._1463_ vssd1 vssd1 vccd1 vccd1 MuI._1464_ sky130_fd_sc_hd__o21a_1
XAuI._1529_ AuI._0711_ AuI._0712_ vssd1 vssd1 vccd1 vccd1 AuI._0713_ sky130_fd_sc_hd__xnor2_1
X_07761_ _00374_ _00376_ _00375_ vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__a21o_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._535_ AuI.pe._045_ AuI.pe._066_ AuI.pe._054_ AuI.pe._056_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._093_ sky130_fd_sc_hd__a22o_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4606_ MuI.b_operand\[20\] MuI._3372_ vssd1 vssd1 vccd1 vccd1 MuI._0310_ sky130_fd_sc_hd__nand2_1
X_09500_ _02124_ _02125_ _02126_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nand3_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06712_ net109 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__buf_2
XMuI._5586_ MuI._3403_ MuI._3397_ MuI._3371_ MuI._0110_ vssd1 vssd1 vccd1 vccd1 MuI._1388_
+ sky130_fd_sc_hd__and4_1
X_07692_ net55 net115 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__nand2_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4028__B MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._466_ AuI.pe._028_ AuI.pe._030_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._031_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4537_ MuI._0103_ MuI._0102_ vssd1 vssd1 vccd1 vccd1 MuI._0234_ sky130_fd_sc_hd__nor2_1
X_09431_ _02046_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__or2b_1
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07930__C _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4970__C MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4468_ MuI.a_operand\[19\] MuI.a_operand\[18\] MuI._2884_ MuI._2880_ vssd1 vssd1
+ vccd1 vccd1 MuI._0158_ sky130_fd_sc_hd__and4_1
X_09362_ _01936_ _01935_ _01928_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4092__A2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6207_ MuI._2067_ MuI._2070_ vssd1 vssd1 vccd1 vccd1 MuI._2071_ sky130_fd_sc_hd__and2_1
XFILLER_178_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07004__A _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _00927_ _00929_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__and2b_1
XMuI._4399_ MuI._2473_ MuI._2374_ vssd1 vssd1 vccd1 vccd1 MuI._0082_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07457__A1 _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _01794_ _01897_ _01896_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a21o_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07457__B2 _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6138_ MuI._1993_ MuI._1909_ MuI._1915_ vssd1 vssd1 vccd1 vccd1 MuI._1995_ sky130_fd_sc_hd__and3_1
XFILLER_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08244_ _00858_ _00861_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__and2_1
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06843__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3883__A MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6069_ MuI._1881_ MuI._1882_ MuI._1918_ vssd1 vssd1 vccd1 vccd1 MuI._1919_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08175_ _00375_ _00376_ _00374_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08406__B1 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07126_ _02020_ _06023_ _02140_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nand3_2
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ _06034_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07674__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10812__B _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4864__D MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13466__B1 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07959_ _00575_ _00576_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__nand2_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ _03527_ _03528_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21o_1
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _02237_ _02265_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__and3_1
XANTENNA__11492__A2 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _05501_ _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5695__D MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _05431_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07999__A2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _04302_ _04303_ _04182_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__o21ai_1
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12992__A2 _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._425__A1 AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._146_ FuI._008_ net152 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[17\] sky130_fd_sc_hd__dlxtn_1
XANTENNA_MuI._3793__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0900_ net60 net28 vssd1 vssd1 vccd1 vccd1 AuI._0120_ sky130_fd_sc_hd__and2b_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ _04226_ _04227_ _04228_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__A _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._077_ FuI._033_ FuI._039_ FuI._042_ vssd1 vssd1 vccd1 vccd1 FuI._043_ sky130_fd_sc_hd__and3b_1
XFILLER_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _00770_ _00800_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__a21oi_2
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._0831_ net109 vssd1 vssd1 vccd1 vccd1 AuI._0051_ sky130_fd_sc_hd__inv_2
X_11384_ _02566_ _02568_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__or2_1
XFILLER_192_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__B1 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _06020_ _06022_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__or2_1
XFILLER_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10335_ _03067_ _01206_ _00445_ _00550_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__nand4_1
XANTENNA__07620__A1 _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07620__B2 _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _05875_ _05876_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__and2b_1
XFILLER_106_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10266_ _00673_ _00710_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__nand2_1
XFILLER_121_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3770_ MuI._0779_ MuI._1021_ MuI._2867_ MuI._2869_ vssd1 vssd1 vccd1 vccd1 MuI._2870_
+ sky130_fd_sc_hd__and4_1
X_12005_ _04823_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10197_ _04262_ _02388_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__or2b_1
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5440_ MuI._1217_ MuI._1225_ MuI._1226_ vssd1 vssd1 vccd1 vccd1 MuI._1227_ sky130_fd_sc_hd__nand3_2
XFILLER_207_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1314_ AuI._0483_ AuI._0510_ AuI._0511_ vssd1 vssd1 vccd1 vccd1 AuI._0512_ sky130_fd_sc_hd__o21a_1
XFILLER_93_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6048__B1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__A _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5371_ MuI._1122_ MuI._1123_ MuI._1138_ vssd1 vssd1 vccd1 vccd1 MuI._1151_ sky130_fd_sc_hd__a21o_1
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08846__C _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _05691_ _05692_ _05792_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__or3_1
XAuI._1245_ AuI._0436_ AuI._0447_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[9\]
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_MuI._6344__A MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4322_ MuI._3418_ MuI._3420_ vssd1 vssd1 vccd1 vccd1 MuI._3422_ sky130_fd_sc_hd__and2b_1
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11272__C _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12838_ _05718_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1176_ AuI._0370_ AuI._0372_ AuI._0375_ AuI._0288_ AuI._0249_ vssd1 vssd1 vccd1
+ vccd1 AuI._0382_ sky130_fd_sc_hd__a221o_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09428__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4253_ MuI._1285_ MuI._2385_ MuI._3352_ MuI._3350_ vssd1 vssd1 vccd1 vccd1 MuI._3353_
+ sky130_fd_sc_hd__a31o_1
XFILLER_203_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _05629_ _05630_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nor3b_1
XANTENNA__08636__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08100__A2 _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4184_ MuI._3283_ MuI._3173_ vssd1 vssd1 vccd1 vccd1 MuI._3284_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10443__B1 _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 a_operand[23] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_6
Xinput31 a_operand[4] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 b_operand[14] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
Xinput53 b_operand[24] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_2
Xinput64 b_operand[5] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_8
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11943__B1 _04604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__D _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09980_ _02041_ _02622_ _02631_ _02644_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a211o_4
XFILLER_131_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4534__B1 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6825_ MuI._2744_ vssd1 vssd1 vccd1 vccd1 MuI.result\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _01518_ _01520_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__and2_1
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6756_ MuI._2654_ vssd1 vssd1 vccd1 vccd1 MuI._2675_ sky130_fd_sc_hd__inv_2
XMuI._3968_ MuI._0350_ MuI._2898_ MuI._2874_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._3068_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _01472_ _01479_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__xor2_1
XANTENNA__11171__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5707_ MuI._2429_ MuI._0327_ MuI._2885_ MuI._3307_ vssd1 vssd1 vccd1 vccd1 MuI._1521_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11171__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _00195_ _00202_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__nand2_1
XMuI._6687_ MuI._3304_ MuI._2598_ vssd1 vssd1 vccd1 vccd1 MuI._2599_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3899_ MuI._1307_ MuI._1802_ MuI._2616_ MuI._2671_ vssd1 vssd1 vccd1 vccd1 MuI._2999_
+ sky130_fd_sc_hd__nand4_1
X_08793_ _01407_ _01409_ _01408_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__o21a_1
XFILLER_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5638_ MuI._1433_ MuI._1434_ MuI._1444_ vssd1 vssd1 vccd1 vccd1 MuI._1445_ sky130_fd_sc_hd__nor3_1
X_07744_ _06452_ _06457_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__nor2_1
XAuI.pe._518_ AuI.pe._077_ vssd1 vssd1 vccd1 vccd1 AuI.pe._078_ sky130_fd_sc_hd__buf_2
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5569_ MuI._1323_ MuI._1324_ MuI._1325_ vssd1 vssd1 vccd1 vccd1 MuI._1369_ sky130_fd_sc_hd__o21bai_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07675_ _00288_ _00291_ _00292_ _06443_ vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__and4bb_1
XFILLER_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._449_ AuI.pe._370_ AuI.pe._374_ AuI.pe._375_ AuI.pe._015_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._016_ sky130_fd_sc_hd__or4_1
X_09414_ _02032_ _02033_ _02024_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__nor3b_2
XANTENNA__10682__B1 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3597__B MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._655__A1 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ _01844_ _01960_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__and2b_1
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12575__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__A _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ _02550_ _04316_ _01892_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a31o_1
XFILLER_194_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ _00819_ _00834_ _00833_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__a21o_1
XFILLER_181_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09884__A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _00773_ _00774_ _00775_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__nand3b_1
XFILLER_162_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07109_ _06418_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[23\] sky130_fd_sc_hd__clkbuf_2
X_08089_ _00705_ _00706_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__or2_2
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__buf_2
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10542__B _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09108__B _01378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6148__B MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5052__B MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06748__A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10945__B_N _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _03651_ _03654_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nand2_2
XFILLER_204_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1030_ net116 net16 net37 net5 AuI._0123_ AuI._0175_ vssd1 vssd1 vccd1 vccd1
+ AuI._0242_ sky130_fd_sc_hd__mux4_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10884_ _03614_ _03616_ _03599_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__a21o_1
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ _02856_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__or2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0812__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07579__A _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12554_ _05039_ _05151_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__or3_1
XFILLER_185_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _04127_ _04270_ _04285_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o211ai_2
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12485_ _05213_ _05215_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and2b_1
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._129_ FuI._010_ net135 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[0\] sky130_fd_sc_hd__dlxtn_1
XANTENNA__12178__B1 _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__D _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11436_ _04211_ _04209_ _04210_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or3_1
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4940_ MuI._0674_ MuI._0676_ vssd1 vssd1 vccd1 vccd1 MuI._0677_ sky130_fd_sc_hd__or2_1
XFILLER_153_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A1 _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09594__B2 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11829__A _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0814_ net51 AuI._0030_ net19 vssd1 vssd1 vccd1 vccd1 AuI._0034_ sky130_fd_sc_hd__or3b_1
X_11367_ _04136_ _04137_ _04096_ _04097_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a211o_1
XFILLER_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4516__B1 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ AuI.result\[23\] _02732_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_
+ sky130_fd_sc_hd__a211o_1
XMuI._4871_ MuI._0425_ MuI._0600_ vssd1 vssd1 vccd1 vccd1 MuI._0601_ sky130_fd_sc_hd__nor2_1
XFILLER_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1362__B AuI._0550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10318_ _02959_ _00421_ _00534_ _00217_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a22o_1
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11298_ _04061_ _04062_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21o_1
XANTENNA__12371__C_N _05218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__A _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6610_ MuI._1814_ MuI._2511_ MuI._1809_ vssd1 vssd1 vccd1 vccd1 MuI._2514_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3822_ MuI._2915_ MuI._2921_ vssd1 vssd1 vccd1 vccd1 MuI._2922_ sky130_fd_sc_hd__xnor2_2
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ net134 _04627_ _03675_ _05467_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__a221o_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _02934_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__buf_2
XFILLER_67_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11267__C _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6541_ MuI._2414_ MuI._2427_ MuI._2437_ vssd1 vssd1 vccd1 vccd1 MuI._2438_ sky130_fd_sc_hd__or3b_1
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3753_ MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 MuI._2853_ sky130_fd_sc_hd__buf_2
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08857__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6472_ MuI._2349_ MuI._2360_ MuI._2361_ vssd1 vssd1 vccd1 vccd1 MuI._2362_ sky130_fd_sc_hd__a21oi_1
XMuI._3684_ MuI._2748_ MuI._2782_ MuI._2781_ vssd1 vssd1 vccd1 vccd1 MuI._2784_ sky130_fd_sc_hd__a21o_1
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5423_ MuI._2869_ MuI._0444_ MuI.a_operand\[1\] MuI._2867_ vssd1 vssd1 vccd1
+ vccd1 MuI._1209_ sky130_fd_sc_hd__a22oi_1
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3698__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5354_ MuI._0085_ MuI._3262_ MuI._0020_ MuI._2341_ vssd1 vssd1 vccd1 vccd1 MuI._1133_
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__12098__C _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1228_ AuI._0398_ AuI._0400_ AuI._0418_ AuI._0431_ vssd1 vssd1 vccd1 vccd1 AuI._0432_
+ sky130_fd_sc_hd__o31a_1
X_07460_ _00077_ _04251_ _00073_ _00075_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08295__D _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4305_ MuI._3269_ MuI._0504_ MuI._3263_ MuI._3404_ vssd1 vssd1 vccd1 vccd1 MuI._3405_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._637__A1 AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._637__B2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5285_ MuI._0928_ MuI._0952_ MuI._1055_ MuI._1056_ vssd1 vssd1 vccd1 vccd1 MuI._1057_
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11208__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1159_ AuI._0364_ AuI._0365_ AuI._0362_ vssd1 vssd1 vccd1 vccd1 AuI._0366_ sky130_fd_sc_hd__a21o_1
X_07391_ _02851_ _04918_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__nand2_1
XFILLER_210_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4236_ MuI._3333_ MuI._3335_ vssd1 vssd1 vccd1 vccd1 MuI._3336_ sky130_fd_sc_hd__and2_1
X_09130_ _03067_ _03917_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__nand2_1
XANTENNA__09282__B1 _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4167_ MuI._3265_ MuI._3266_ vssd1 vssd1 vccd1 vccd1 MuI._3267_ sky130_fd_sc_hd__xor2_1
X_09061_ _01677_ _01678_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__nor2_1
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07639__D _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08012_ _00531_ _00532_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__nor2_1
XMuI._4098_ MuI._2671_ MuI._2841_ vssd1 vssd1 vccd1 vccd1 MuI._3198_ sky130_fd_sc_hd__nand2_1
XFILLER_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09034__B1 _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__A1 _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__B2 _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ _02603_ _02597_ _02609_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__or3_1
XFILLER_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07655__C _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6808_ MuI._0141_ MuI._2502_ MuI._0130_ vssd1 vssd1 vccd1 vccd1 MuI._2732_ sky130_fd_sc_hd__a21oi_2
X_08914_ _01508_ _01509_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__and4bb_1
XANTENNA__13133__A2 _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ _02516_ _02526_ _02552_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o21ai_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__B1 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6739_ MuI._2643_ MuI._2647_ MuI._2655_ vssd1 vssd1 vccd1 vccd1 MuI._2656_ sky130_fd_sc_hd__and3_1
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07952__A _00567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _06548_ _04832_ _04896_ _02291_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a22oi_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11474__A _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08776_ _03024_ _04057_ _01385_ _01384_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__a31o_2
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07727_ net55 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__buf_4
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07658_ _00261_ _00264_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4216__B MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._628__A1 AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07589_ _00204_ _00205_ _00206_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__nand3_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09328_ _01939_ _01943_ _01944_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a211oi_4
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08076__A1 _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08076__B2 _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09259_ _01875_ _01874_ _01672_ _01665_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a211o_1
XFILLER_194_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08007__B _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12270_ _05107_ _05108_ _04970_ _04973_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a211o_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _03979_ _03959_ _03961_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__and3_1
XFILLER_181_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07846__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09119__A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _03632_ _03807_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__or2_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _05402_ _03293_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__and2b_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11083_ _03830_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__nor2_1
XFILLER_89_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3721__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A a_operand[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3721__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5998__A MuI._1836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _00816_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__xor2_2
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12883__A1 _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__A2 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0807__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__A2 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12635__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ _04784_ _04785_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3949__C MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__B2 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ _04197_ _02941_ _02731_ AuI.result\[4\] vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12927__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._1013_ AuI._0199_ AuI._0200_ AuI._0224_ AuI._0176_ vssd1 vssd1 vccd1 vccd1 AuI._0225_
+ sky130_fd_sc_hd__a31oi_1
XFILLER_182_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _03447_ _03457_ _03456_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10728__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5070_ MuI._2838_ MuI._0304_ MuI._0444_ MuI._2836_ vssd1 vssd1 vccd1 vccd1 MuI._0820_
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12646__C _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09301__B _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12606_ _05469_ _05470_ _05333_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__a21oi_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1357__B AuI._0550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__A1 _02815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4021_ MuI._3088_ MuI._3089_ MuI._3119_ MuI._3120_ vssd1 vssd1 vccd1 vccd1 MuI._3121_
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _06439_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__buf_2
XFILLER_157_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07102__A _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _03489_ _05389_ _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a21o_1
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11610__A2 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12468_ _05320_ _05321_ _05191_ _05195_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__o211ai_2
XANTENNA__06941__A _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12662__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5972_ MuI._1795_ MuI._1810_ MuI._1811_ vssd1 vssd1 vccd1 vccd1 MuI._1812_ sky130_fd_sc_hd__a21o_1
X_11419_ _04191_ _04192_ _04188_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21o_1
XFILLER_125_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07756__B _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12399_ _02800_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__inv_2
XFILLER_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4923_ MuI._0649_ MuI._0651_ MuI._0657_ vssd1 vssd1 vccd1 vccd1 MuI._0659_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10182__B _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._783_ AuI.pe._016_ AuI.pe._299_ vssd1 vssd1 vccd1 vccd1 AuI.pe._324_ sky130_fd_sc_hd__nand2_1
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4854_ MuI._0580_ MuI._0582_ vssd1 vssd1 vccd1 vccd1 MuI._0583_ sky130_fd_sc_hd__and2_1
XFILLER_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06960_ _04994_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__and3_1
XFILLER_140_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3805_ MuI._2888_ MuI._2897_ MuI._2903_ vssd1 vssd1 vccd1 vccd1 MuI._2905_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4785_ MuI._0503_ MuI._0506_ vssd1 vssd1 vccd1 vccd1 MuI._0507_ sky130_fd_sc_hd__nor2_1
XFILLER_67_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06891_ _04251_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6524_ MuI._2209_ MuI._2275_ vssd1 vssd1 vccd1 vccd1 MuI._2420_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3736_ MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 MuI._2836_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11294__A _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _01246_ _01247_ _06608_ _04369_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__and4bb_1
XFILLER_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07491__B net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4268__A2 MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6455_ MuI._1948_ MuI._1947_ vssd1 vssd1 vccd1 vccd1 MuI._2344_ sky130_fd_sc_hd__and2b_1
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3667_ MuI.b_operand\[13\] vssd1 vssd1 vccd1 vccd1 MuI._2693_ sky130_fd_sc_hd__buf_2
X_08561_ _01175_ _01177_ _01178_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__nor3_1
XFILLER_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5406_ MuI._2895_ MuI._3372_ vssd1 vssd1 vccd1 vccd1 MuI._1190_ sky130_fd_sc_hd__nand2_1
X_07512_ _00086_ _00081_ _00047_ _04638_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__and4_1
XMuI._6386_ MuI._1887_ MuI._2851_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._2268_ sky130_fd_sc_hd__nand3b_1
XFILLER_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3598_ MuI._0746_ MuI._0801_ MuI._1164_ MuI._0581_ vssd1 vssd1 vccd1 vccd1 MuI._1934_
+ sky130_fd_sc_hd__a22oi_1
X_08492_ _00926_ _00925_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__and2b_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4036__B MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12837__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5337_ MuI._0978_ MuI._0980_ vssd1 vssd1 vccd1 vccd1 MuI._1114_ sky130_fd_sc_hd__nor2_1
XANTENNA_AuI.pe._404__A AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07443_ _02894_ _02948_ _04703_ _04778_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__and4_1
XFILLER_90_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5268_ MuI._2429_ MuI.b_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._1038_ sky130_fd_sc_hd__nand2_1
XFILLER_149_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ _06659_ _06660_ _06673_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__and3_1
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4219_ MuI._3316_ MuI._3317_ MuI._3318_ vssd1 vssd1 vccd1 vccd1 MuI._3319_ sky130_fd_sc_hd__o21ba_1
X_09113_ _01710_ _01709_ _01708_ _01696_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__o211a_1
XANTENNA__07012__A net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5199_ MuI._2895_ MuI._3363_ MuI._0796_ MuI._0797_ vssd1 vssd1 vccd1 vccd1 MuI._0962_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3594__C MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09044_ _01659_ _01660_ _01646_ _01585_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a211o_1
XFILLER_191_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06851__A _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13354__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07385__C _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13106__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09946_ _02592_ _02605_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__or2_2
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08778__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _02531_ _02533_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__nor2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1385__A2 AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _01438_ _01440_ _01439_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o21ai_1
XANTENNA_MuI._5456__A1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5456__B2 MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09652__A2_N _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08759_ _01375_ _01376_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__nor2_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ _04405_ _04415_ _04414_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a21o_1
XFILLER_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10170__B_N _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07656__A1_N _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _02388_ _05895_ _05970_ _02345_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11651__B _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10548__A _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _03842_ _05917_ _06322_ _06321_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a31o_1
XANTENNA__09121__B _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ _03356_ _03366_ _03367_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and3_1
XFILLER_139_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6161__B MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5058__A MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1427__A_N AuI._0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ _06281_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xor2_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _00816_ _03124_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__and2b_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08960__B _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12322_ _05164_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nor2_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06761__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _05090_ _05091_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__xor2_4
XFILLER_170_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3942__A1 MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _01147_ _01146_ _04972_ _05036_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3942__B2 MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1631_ AuI.pe.Significand\[20\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0797_
+ sky130_fd_sc_hd__or2_1
XFILLER_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5505__B MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ _02845_ _04898_ _02846_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI._1073__A1 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _03882_ _03886_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nand3_2
XAuI._1562_ AuI._0606_ AuI._0739_ AuI._0740_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[7\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0820__B2 net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11066_ _03776_ _03778_ _03812_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1493_ AuI._0375_ AuI._0498_ AuI._0577_ vssd1 vssd1 vccd1 vccd1 AuI._0679_ sky130_fd_sc_hd__or3b_1
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4570_ MuI._0267_ MuI._0269_ vssd1 vssd1 vccd1 vccd1 MuI._0270_ sky130_fd_sc_hd__xnor2_1
X_10017_ _02674_ _02684_ _01878_ _01876_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__o211a_1
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3521_ MuI._1065_ MuI._1054_ vssd1 vssd1 vccd1 vccd1 MuI._1087_ sky130_fd_sc_hd__and2b_1
XFILLER_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4782__D MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4137__A MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6240_ MuI._2102_ MuI._2103_ MuI._2106_ vssd1 vssd1 vccd1 vccd1 MuI._2107_ sky130_fd_sc_hd__nand3_1
XMuI._3452_ MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 MuI._0328_ sky130_fd_sc_hd__buf_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06936__A _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _04781_ _04782_ _04783_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a21o_1
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12657__B _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6171_ MuI._2028_ MuI._2029_ MuI._2030_ vssd1 vssd1 vccd1 vccd1 MuI._2031_ sky130_fd_sc_hd__o21bai_1
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _03651_ _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__xor2_4
X_11899_ _04709_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__xor2_1
XMuI._5122_ MuI._0874_ MuI._0875_ MuI._0873_ vssd1 vssd1 vccd1 vccd1 MuI._0877_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10177__B _02848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5053_ MuI._3189_ MuI._3190_ MuI.a_operand\[6\] MuI.a_operand\[5\] vssd1 vssd1
+ vccd1 vccd1 MuI._0802_ sky130_fd_sc_hd__and4_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4004_ MuI._3100_ MuI._3101_ MuI._3102_ vssd1 vssd1 vccd1 vccd1 MuI._3104_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07767__A net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ _06377_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_117_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11347__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11347__B2 _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5955_ MuI._1770_ MuI._1793_ vssd1 vssd1 vccd1 vccd1 MuI._1794_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._4957__D MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__B_N _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4906_ MuI._2814_ MuI._2813_ MuI._0111_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._0640_
+ sky130_fd_sc_hd__and4_1
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _02422_ _02413_ _02421_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nand3_1
XMuI._5886_ MuI._1660_ MuI._1662_ vssd1 vssd1 vccd1 vccd1 MuI._1718_ sky130_fd_sc_hd__nor2_1
XFILLER_114_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07992_ _00607_ _00608_ _00609_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a21o_1
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._766_ AuI.pe._105_ AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 AuI.pe._310_ sky130_fd_sc_hd__or2_1
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4837_ MuI._2852_ MuI.a_operand\[15\] MuI._2884_ MuI._2880_ vssd1 vssd1 vccd1
+ vccd1 MuI._0564_ sky130_fd_sc_hd__and4_1
X_06943_ _04811_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[13\] sky130_fd_sc_hd__clkbuf_1
X_09731_ _02366_ _02374_ _02307_ _02375_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__o211a_2
XANTENNA__11736__B _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10307__C1 _00702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._697_ AuI.pe._089_ AuI.pe._150_ AuI.pe._173_ AuI.pe._062_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._244_ sky130_fd_sc_hd__a22o_1
XFILLER_83_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4768_ MuI._0286_ MuI._0487_ vssd1 vssd1 vccd1 vccd1 MuI._0488_ sky130_fd_sc_hd__xnor2_1
X_09662_ _02293_ _02300_ _02301_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a21bo_1
X_06874_ _04068_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__and3_1
XANTENNA__08748__D _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__C _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6507_ MuI._2211_ MuI._2212_ vssd1 vssd1 vccd1 vccd1 MuI._2401_ sky130_fd_sc_hd__nor2_1
XFILLER_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3719_ MuI._2816_ MuI._2818_ vssd1 vssd1 vccd1 vccd1 MuI._2819_ sky130_fd_sc_hd__nor2_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08613_ _01229_ _01230_ _02712_ _04585_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__and4bb_1
XANTENNA__07007__A _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4699_ MuI._0409_ MuI._0410_ MuI._0411_ vssd1 vssd1 vccd1 vccd1 MuI._0412_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09593_ _06513_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__buf_4
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6438_ MuI._2258_ MuI._2261_ MuI._2259_ vssd1 vssd1 vccd1 vccd1 MuI._2325_ sky130_fd_sc_hd__o21ba_1
XFILLER_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _00262_ _00303_ _01099_ _01100_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6369_ MuI._2247_ MuI._2248_ vssd1 vssd1 vccd1 vccd1 MuI._2249_ sky130_fd_sc_hd__or2_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08475_ _01077_ _01078_ _01090_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11822__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _00037_ _00042_ _00043_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__or3_1
XANTENNA__08483__D _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09779__A1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B1 _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10518__D _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ _06649_ _06650_ _06655_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a21o_1
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0910__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__A1 _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11586__B2 _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__C _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07288_ _06578_ _06579_ _06581_ _05101_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__and4_1
XFILLER_191_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09027_ _01643_ _01642_ _01627_ _01547_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a211oi_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12535__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11927__A _04721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__A1_N _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4986__A2_N MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ _02328_ _02588_ _02589_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__nand3_1
XFILLER_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11646__B _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10550__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12940_ _05779_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__xnor2_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _02630_ _02622_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12758__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ MuI.result\[10\] _02737_ _04011_ _02860_ _04628_ vssd1 vssd1 vccd1 vccd1
+ _04629_ sky130_fd_sc_hd__a221o_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06756__A _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3796__A MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11753_ _04551_ _04552_ _04499_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _06461_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__clkbuf_4
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _04477_ _04479_ _04298_ _04363_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__a211oi_4
XANTENNA__07493__A2 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13423_ _02817_ _02915_ _02919_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o21bai_2
X_10635_ _03348_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__xor2_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._470__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _03561_ _02724_ _06262_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__a211o_1
XANTENNA__08907__A1_N _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10566_ _03219_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__xor2_1
XANTENNA_AuI._1294__A1 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0993_ AuI._0143_ AuI._0204_ vssd1 vssd1 vccd1 vccd1 AuI._0205_ sky130_fd_sc_hd__and2_2
X_12305_ _05050_ _05048_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__or2b_1
XFILLER_127_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13318__A2 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13285_ _06166_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__xor2_1
X_10497_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10444__C _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12236_ _05071_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__xor2_1
XFILLER_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5740_ MuI._0990_ MuI._1551_ MuI._1550_ vssd1 vssd1 vccd1 vccd1 MuI._1557_ sky130_fd_sc_hd__a21bo_1
XFILLER_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1614_ AuI.pe.Significand\[16\] AuI._0695_ AuI._0760_ AuI._0783_ vssd1 vssd1
+ vccd1 vccd1 AuI.result\[16\] sky130_fd_sc_hd__o211a_1
X_12167_ _04999_ _04880_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__and2b_1
XAuI.pe._620_ AuI.pe.significand\[10\] AuI.pe._149_ AuI.pe._395_ AuI.pe._105_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._172_ sky130_fd_sc_hd__and4b_1
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5671_ MuI._1002_ MuI._1007_ vssd1 vssd1 vccd1 vccd1 MuI._1481_ sky130_fd_sc_hd__and2_1
X_11118_ _03867_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__xor2_4
XANTENNA_MuI._3679__B1 MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1545_ AuI._0606_ AuI._0725_ AuI._0726_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[4\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12098_ _00921_ _01206_ _05649_ _03449_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nand4_1
XANTENNA__08211__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._551_ AuI.pe._106_ AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 AuI.pe._108_ sky130_fd_sc_hd__nand2_1
XANTENNA__10460__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4622_ MuI.a_operand\[12\] vssd1 vssd1 vccd1 vccd1 MuI._0327_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._5251__A MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11049_ _03792_ _03793_ _03785_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a21o_1
XFILLER_49_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1476_ AuI._0415_ AuI._0411_ vssd1 vssd1 vccd1 vccd1 AuI._0662_ sky130_fd_sc_hd__or2b_1
Xinput7 a_operand[11] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_8
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07705__B1 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4891__A2 MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._482_ AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 AuI.pe._045_ sky130_fd_sc_hd__buf_2
XFILLER_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4553_ MuI._0249_ MuI._0250_ vssd1 vssd1 vccd1 vccd1 MuI._0252_ sky130_fd_sc_hd__or2_1
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09170__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07181__A1 _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3504_ MuI._0757_ MuI._0856_ MuI._0889_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._0900_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07181__B2 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4484_ MuI._0158_ MuI._0160_ MuI._0175_ vssd1 vssd1 vccd1 vccd1 MuI._0176_ sky130_fd_sc_hd__o21ai_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6223_ MuI._1142_ MuI._2916_ MuI._2627_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._2089_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12387__B _05233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3435_ MuI._0119_ MuI._0130_ vssd1 vssd1 vccd1 vccd1 MuI._0141_ sky130_fd_sc_hd__nor2_1
XFILLER_205_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6154_ MuI._1032_ MuI._2473_ vssd1 vssd1 vccd1 vccd1 MuI._2013_ sky130_fd_sc_hd__nand2_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _06599_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__buf_4
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08881__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5105_ MuI._2374_ MuI._2895_ vssd1 vssd1 vccd1 vccd1 MuI._0859_ sky130_fd_sc_hd__nand2_1
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07211_ _06485_ _06510_ _06509_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__a21o_1
XMuI._6085_ MuI._1930_ MuI._1936_ vssd1 vssd1 vccd1 vccd1 MuI._1937_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08191_ _00807_ _00808_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__xnor2_2
XANTENNA_MuI._6810__A MuI._2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5036_ MuI._0671_ MuI._0666_ MuI._0670_ vssd1 vssd1 vccd1 vccd1 MuI._0783_ sky130_fd_sc_hd__nand3_1
XANTENNA__11568__B2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ _04035_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__buf_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__C _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07073_ _06202_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10354__C _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5938_ MuI._1743_ MuI._1744_ MuI._1745_ vssd1 vssd1 vccd1 vccd1 MuI._1775_ sky130_fd_sc_hd__a21oi_1
XFILLER_102_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._818_ AuI.pe._345_ AuI.pe._348_ AuI.pe._350_ AuI.pe._356_ AuI.operand_a\[26\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._357_ sky130_fd_sc_hd__a41o_1
XANTENNA__07944__B1 _00105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5869_ MuI._1696_ MuI._1697_ MuI._1622_ MuI._1684_ vssd1 vssd1 vccd1 vccd1 MuI._1699_
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ net118 net117 _00592_ _00089_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__and4_1
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._749_ AuI.pe.significand\[22\] AuI.pe._291_ vssd1 vssd1 vccd1 vccd1 AuI.pe._293_
+ sky130_fd_sc_hd__nor2_1
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _06460_ _04165_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__and2_1
X_06926_ net7 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__buf_4
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12296__A2 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _02277_ _02282_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a21oi_1
X_06857_ _03884_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__buf_4
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11482__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4208__C MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ _02120_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a21oi_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__C _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ net49 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__buf_4
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08527_ _01144_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10098__A _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._799__A AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _00886_ _01069_ _01068_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__a21o_1
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07409_ _00025_ _00024_ _06641_ _06576_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__o211ai_2
XFILLER_196_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10248__D _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08389_ _01004_ _01005_ _01006_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__nand3_2
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._093_ FuI.a_operand\[27\] FuI.a_operand\[28\] FuI.a_operand\[29\] net105 vssd1
+ vssd1 vccd1 vccd1 FuI._054_ sky130_fd_sc_hd__or4b_2
X_10420_ _00810_ _00811_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__nor2_1
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07227__A2 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5347__B1 MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07200__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ _06610_ _05198_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nand2_1
XFILLER_137_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12508__B1 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13070_ _05891_ _05892_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__o21ai_1
X_10282_ _06429_ _04122_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI._1028__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12021_ _04839_ _04840_ _04841_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__a21o_1
XANTENNA__08727__A2 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07573__C _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5071__A MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1330_ AuI._0518_ AuI._0524_ AuI._0525_ AuI._0257_ vssd1 vssd1 vccd1 vccd1 AuI._0526_
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__A2 _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13484__B2 _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12923_ _03744_ _05456_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__nand3_1
XAuI._1261_ AuI._0438_ AuI._0335_ AuI._0421_ AuI._0461_ vssd1 vssd1 vccd1 vccd1 AuI._0462_
+ sky130_fd_sc_hd__o211a_2
XFILLER_207_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07163__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07163__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4118__C MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1192_ AuI._0396_ AuI._0397_ vssd1 vssd1 vccd1 vccd1 AuI._0398_ sky130_fd_sc_hd__nand2b_2
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12854_ _05648_ _05651_ _05736_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or3_1
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13236__B2 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _04606_ _04609_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__or2_1
XANTENNA_output100_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__B _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _05661_ _05662_ _05599_ _05600_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o211a_1
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11736_ _00088_ _05380_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__nand2_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _04278_ _04282_ _04460_ _04461_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__a211o_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13406_ _02917_ _02875_ _06108_ _06228_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__o22a_1
X_10618_ _03135_ _03289_ _03330_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a21oi_2
X_11598_ _00046_ _03424_ _03425_ _00049_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a22o_1
XFILLER_183_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10455__B _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07110__A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10549_ _06545_ _03257_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__nand2_1
X_13337_ _03842_ _05724_ _06182_ _06179_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__a31o_1
XAuI._0976_ AuI._0185_ AuI._0187_ AuI._0175_ vssd1 vssd1 vccd1 vccd1 AuI._0188_ sky130_fd_sc_hd__mux2_1
XFILLER_109_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6841_ MuI._2680_ MuI._2684_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI.result\[13\]
+ sky130_fd_sc_hd__nor3b_1
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6776__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13268_ _03755_ _05777_ _06175_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__a21o_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6772_ MuI._2691_ MuI._2689_ MuI._2621_ MuI._2683_ vssd1 vssd1 vccd1 vccd1 MuI._2692_
+ sky130_fd_sc_hd__a2bb2o_1
XMuI._3984_ MuI._3082_ MuI._3083_ vssd1 vssd1 vccd1 vccd1 MuI._3084_ sky130_fd_sc_hd__or2_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__nor2_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13199_ _05947_ _06041_ _06104_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5723_ MuI._1518_ MuI._1536_ MuI._1537_ vssd1 vssd1 vccd1 vccd1 MuI._1539_ sky130_fd_sc_hd__and3_1
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._603_ AuI.pe._037_ AuI.pe._146_ AuI.pe._148_ AuI.pe._156_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[12\] sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11717__D _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5654_ MuI._0984_ MuI._1060_ vssd1 vssd1 vccd1 vccd1 MuI._1463_ sky130_fd_sc_hd__nand2_1
XAuI._1528_ AuI._0655_ AuI._0652_ vssd1 vssd1 vccd1 vccd1 AuI._0712_ sky130_fd_sc_hd__and2b_1
X_07760_ _00152_ _00154_ _00151_ vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__o21bai_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5412__C MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._534_ AuI.pe._074_ AuI.pe._085_ AuI.pe._088_ AuI.pe._092_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[7\] sky130_fd_sc_hd__o22a_1
XFILLER_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4605_ MuI._0867_ MuI._0111_ MuI._0308_ vssd1 vssd1 vccd1 vccd1 MuI._0309_ sky130_fd_sc_hd__and3_1
XFILLER_110_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4309__B MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _02313_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[3\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07780__A _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5585_ MuI._3397_ MuI._0305_ MuI._0111_ MuI._3403_ vssd1 vssd1 vccd1 vccd1 MuI._1387_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07691_ _00278_ _03432_ net132 _06430_ vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__and4_1
XAuI._1459_ AuI._0411_ AuI._0415_ vssd1 vssd1 vccd1 vccd1 AuI._0645_ sky130_fd_sc_hd__or2b_1
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._465_ AuI.pe._014_ vssd1 vssd1 vccd1 vccd1 AuI.pe._030_ sky130_fd_sc_hd__buf_2
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4536_ MuI._2817_ MuI._3372_ MuI._0232_ vssd1 vssd1 vccd1 vccd1 MuI._0233_ sky130_fd_sc_hd__and3_1
X_09430_ _02047_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07930__D _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4467_ MuI._1461_ MuI._2885_ MuI._2881_ MuI.a_operand\[19\] vssd1 vssd1 vccd1
+ vccd1 MuI._0157_ sky130_fd_sc_hd__a22oi_1
X_09361_ _01970_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a21bo_1
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07425__A1_N _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6206_ MuI._2012_ MuI._2069_ vssd1 vssd1 vccd1 vccd1 MuI._2070_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08312_ _00927_ _00929_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__xnor2_1
XMuI._4398_ MuI._0078_ MuI._0079_ MuI._0080_ vssd1 vssd1 vccd1 vccd1 MuI._0081_ sky130_fd_sc_hd__o21ba_1
X_09292_ _01907_ _01909_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__and2_1
XANTENNA__07457__A2 _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6137_ MuI._1909_ MuI._1915_ MuI._1993_ vssd1 vssd1 vccd1 vccd1 MuI._1994_ sky130_fd_sc_hd__a21oi_1
XFILLER_193_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10461__A1 _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _00859_ _00860_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__xnor2_2
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10646__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6068_ MuI._1850_ MuI._1880_ vssd1 vssd1 vccd1 vccd1 MuI._1918_ sky130_fd_sc_hd__and2_1
XFILLER_118_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12564__C _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3883__B MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08174_ _00790_ _00791_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__or2_1
XANTENNA__08406__A1 _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08406__B2 _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5019_ MuI._0589_ MuI._0590_ MuI._0609_ MuI._0610_ vssd1 vssd1 vccd1 vccd1 MuI._0764_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07020__A _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ _06426_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07056_ _06023_ _02140_ _02020_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and3b_1
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10812__C _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4304__A1 MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07958_ _00567_ _00569_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__xor2_1
XFILLER_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06909_ _04445_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__buf_6
XFILLER_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07889_ _03604_ _06433_ _00272_ _00506_ vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22oi_1
XFILLER_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _02214_ _02264_ _02258_ _02263_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__o211ai_1
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09559_ _02172_ _02171_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__and2b_1
XFILLER_197_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._673__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ _03722_ _05209_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__and2_1
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _04182_ _04302_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__or3_1
XFILLER_184_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._145_ FuI._007_ net151 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[16\] sky130_fd_sc_hd__dlxtn_1
XFILLER_7_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3793__B MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11452_ _04226_ _04227_ _04228_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__and3_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10275__B _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._076_ net104 FuI.a_operand\[23\] FuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1
+ FuI._042_ sky130_fd_sc_hd__a21o_1
X_10403_ _00798_ _00799_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._5066__A MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0830_ net108 vssd1 vssd1 vccd1 vccd1 AuI._0050_ sky130_fd_sc_hd__inv_2
XFILLER_165_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11383_ _04154_ _04155_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__or2_1
XFILLER_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__A1 _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A b_operand[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _01206_ _04843_ _04907_ _00921_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__a22o_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__B2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ _06020_ _06022_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__nand2_1
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07620__A2 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _05947_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__and2_1
XFILLER_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10291__A _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _03820_ _04004_ _00689_ _00687_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__a31o_1
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12901__B1 _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _03722_ _04854_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__and2_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5513__B MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _04671_ _02723_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__or2b_1
XFILLER_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1313_ AuI._0484_ AuI._0494_ AuI._0495_ vssd1 vssd1 vccd1 vccd1 AuI._0511_ sky130_fd_sc_hd__o21bai_1
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6048__A1 MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6048__B2 MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5370_ MuI._1145_ MuI._1149_ vssd1 vssd1 vccd1 vccd1 MuI._1150_ sky130_fd_sc_hd__xnor2_1
X_12906_ _05691_ _05692_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__o21ai_1
XAuI._1244_ AuI._0445_ AuI._0446_ vssd1 vssd1 vccd1 vccd1 AuI._0447_ sky130_fd_sc_hd__and2b_1
XFILLER_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08846__D _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6344__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4321_ MuI._3418_ MuI._3420_ vssd1 vssd1 vccd1 vccd1 MuI._3421_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0932__B1 net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1175_ AuI._0366_ AuI._0381_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[5\]
+ sky130_fd_sc_hd__xnor2_4
X_12837_ _03658_ _05456_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__nand2_1
XFILLER_188_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11272__D _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4252_ MuI._3350_ MuI._3351_ vssd1 vssd1 vccd1 vccd1 MuI._3352_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._6063__C MuI._1908_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08636__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06944__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _05643_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08636__B2 _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4183_ MuI._3160_ MuI._3171_ vssd1 vssd1 vccd1 vccd1 MuI._3283_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__A1 _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11719_ _00221_ _05585_ _04514_ _04515_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__nand4_1
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11640__B1 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12699_ _05567_ _05569_ _03133_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__o21a_1
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput10 a_operand[14] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_6
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 a_operand[24] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_4
XFILLER_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10185__B _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput32 a_operand[5] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_2
Xinput43 b_operand[15] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_4
Xinput54 b_operand[25] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_6
XFILLER_190_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput65 b_operand[6] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_2
XFILLER_171_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10109__A_N _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0959_ AuI._0164_ AuI._0169_ AuI._0170_ vssd1 vssd1 vccd1 vccd1 AuI._0171_ sky130_fd_sc_hd__and3_1
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4534__A1 MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6824_ MuI._2685_ MuI._2703_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2744_ sky130_fd_sc_hd__and3_1
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4534__B2 MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08930_ _01546_ _01545_ _01533_ _01495_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__o211a_1
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6755_ MuI._2666_ MuI._2673_ vssd1 vssd1 vccd1 vccd1 MuI._2674_ sky130_fd_sc_hd__or2_1
XMuI._3967_ MuI._2898_ MuI._0515_ MuI._3056_ vssd1 vssd1 vccd1 vccd1 MuI._3067_ sky130_fd_sc_hd__and3_1
X_08861_ _01473_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._6287__A1 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5706_ MuI._2451_ MuI._2892_ MuI._3185_ MuI._2440_ vssd1 vssd1 vccd1 vccd1 MuI._1520_
+ sky130_fd_sc_hd__a22oi_2
XANTENNA_MuI._6287__B2 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11171__A2 _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6686_ MuI._0013_ MuI._2592_ MuI._0791_ vssd1 vssd1 vccd1 vccd1 MuI._2598_ sky130_fd_sc_hd__a21bo_1
X_07812_ _00410_ _00428_ _00429_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4298__B1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3898_ MuI._1263_ MuI._2528_ vssd1 vssd1 vccd1 vccd1 MuI._2998_ sky130_fd_sc_hd__nand2_1
X_08792_ _01407_ _01408_ _01409_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__nor3_1
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5637_ MuI._1413_ MuI._1436_ MuI._1443_ vssd1 vssd1 vccd1 vccd1 MuI._1444_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI.pe._407__A AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _00341_ _00333_ _00359_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__nor3_1
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._517_ AuI.pe.significand\[17\] AuI.pe._000_ AuI.pe._383_ AuI.pe._076_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._077_ sky130_fd_sc_hd__and4_1
XFILLER_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5568_ MuI._1323_ MuI._1324_ MuI._1325_ vssd1 vssd1 vccd1 vccd1 MuI._1368_ sky130_fd_sc_hd__or3b_1
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07674_ net55 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__buf_4
XAuI.pe._448_ AuI.pe._013_ AuI.pe.significand\[2\] AuI.pe.significand\[3\] AuI.pe._014_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._015_ sky130_fd_sc_hd__or4b_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0923__A0 net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4519_ MuI._1263_ MuI._3363_ MuI._0087_ MuI._0089_ vssd1 vssd1 vccd1 vccd1 MuI._0214_
+ sky130_fd_sc_hd__o2bb2a_1
X_09413_ _02030_ _02029_ _02028_ _02021_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__o211a_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10682__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07015__A _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5499_ MuI._1276_ MuI._1282_ MuI._1283_ vssd1 vssd1 vccd1 vccd1 MuI._1292_ sky130_fd_sc_hd__and3_1
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3597__C MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10682__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09344_ _01767_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__xnor2_2
XFILLER_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12575__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08772__C _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _01890_ _01891_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__nor2_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08226_ _00839_ _00843_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _06516_ _06461_ _05638_ _06520_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__a22o_1
XFILLER_181_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09884__B _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07108_ _05467_ _06414_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__and2_1
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07685__A _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _00703_ _00704_ _00491_ _00493_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__o211a_1
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ _05842_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_161_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _02705_ _02720_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__nor2_4
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6148__C MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4828__A2 MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13439__B2 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ _03657_ _03667_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nand2_1
XFILLER_84_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _03599_ _03614_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__nand3_2
XFILLER_204_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08963__B _01407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _05487_ _02901_ _02928_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__mux2_1
XFILLER_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06764__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0812__B net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _05405_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__xor2_1
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11504_ _04283_ _04284_ _04121_ _04126_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__o211ai_1
XFILLER_200_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _05337_ _05339_ _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__o211ai_4
XFILLER_185_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._128_ FuI._032_ vssd1 vssd1 vccd1 vccd1 FuI._013_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12178__A1 _00555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12178__B2 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ _04209_ _04210_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0813_ net50 AuI._0026_ AuI._0031_ AuI._0032_ vssd1 vssd1 vccd1 vccd1 AuI._0033_
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__A2 _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _04096_ _04097_ _04136_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__o211ai_4
XFILLER_153_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4870_ MuI._2583_ MuI._2330_ MuI._0423_ MuI._0424_ vssd1 vssd1 vccd1 vccd1 MuI._0600_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13105_ _05531_ _03675_ _02722_ _03346_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__a22o_1
X_10317_ _00751_ _00754_ _00752_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__o21bai_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11297_ _03950_ _03952_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__nand2_1
XMuI._3821_ MuI._2917_ MuI._2920_ vssd1 vssd1 vccd1 vccd1 MuI._2921_ sky130_fd_sc_hd__and2b_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__B _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ MuI.result\[22\] _02737_ _02707_ _02908_ _05932_ vssd1 vssd1 vccd1 vccd1
+ _05933_ sky130_fd_sc_hd__a221o_1
X_10248_ _06023_ _02020_ _02064_ _02705_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__and4b_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._582__B2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__D _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6540_ MuI._2434_ MuI._2436_ vssd1 vssd1 vccd1 vccd1 MuI._2437_ sky130_fd_sc_hd__and2_1
XMuI._3752_ MuI.a_operand\[16\] vssd1 vssd1 vccd1 vccd1 MuI._2852_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11845__A _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ _02669_ _04607_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__or2b_1
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6471_ MuI._2359_ MuI._2351_ vssd1 vssd1 vccd1 vccd1 MuI._2361_ sky130_fd_sc_hd__and2b_1
XFILLER_120_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3683_ MuI._2748_ MuI._2781_ MuI._2782_ vssd1 vssd1 vccd1 vccd1 MuI._2783_ sky130_fd_sc_hd__nand3_1
XANTENNA__09315__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__C net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5422_ MuI._2871_ MuI.a_operand\[0\] vssd1 vssd1 vccd1 vccd1 MuI._1207_ sky130_fd_sc_hd__nand2_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3698__B MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5353_ MuI._3362_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._1132_ sky130_fd_sc_hd__nand2_1
XFILLER_35_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12098__D _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1227_ AuI._0398_ AuI._0402_ AuI._0418_ AuI._0430_ AuI._0417_ vssd1 vssd1 vccd1
+ vccd1 AuI._0431_ sky130_fd_sc_hd__o32a_1
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4304_ MuI._0339_ MuI._3269_ MuI._3403_ MuI._0504_ vssd1 vssd1 vccd1 vccd1 MuI._3404_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_50_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5284_ MuI._1014_ MuI._1015_ MuI._1052_ MuI._1053_ vssd1 vssd1 vccd1 vccd1 MuI._1056_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1158_ AuI._0364_ AuI._0365_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[4\]
+ sky130_fd_sc_hd__xor2_4
X_07390_ _00004_ _00005_ _00006_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a21o_1
XFILLER_62_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4235_ MuI._3216_ MuI._3334_ vssd1 vssd1 vccd1 vccd1 MuI._3335_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6090__A MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1089_ AuI._0139_ AuI._0298_ AuI._0299_ vssd1 vssd1 vccd1 vccd1 AuI._0300_ sky130_fd_sc_hd__or3b_1
XANTENNA__10196__A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09282__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09282__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4166_ MuI._0790_ MuI._2967_ vssd1 vssd1 vccd1 vccd1 MuI._3266_ sky130_fd_sc_hd__nand2_1
XFILLER_187_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09060_ _01625_ _01622_ _01624_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4322__B MuI._3420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__B_N _00665_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08011_ _00623_ _00624_ _00628_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__a21o_1
XMuI._4097_ MuI._2864_ MuI._3182_ MuI._3196_ vssd1 vssd1 vccd1 vccd1 MuI._3197_ sky130_fd_sc_hd__a21o_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09034__A1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09034__B2 _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09585__A2 _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _02585_ _02625_ _02597_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__or3_1
XFILLER_171_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07655__D _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6807_ MuI._2672_ MuI._2674_ MuI._2730_ vssd1 vssd1 vccd1 vccd1 MuI._2731_ sky130_fd_sc_hd__and3_1
X_08913_ _01528_ _01529_ _01510_ _01511_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a211o_1
XMuI._4999_ MuI.a_operand\[16\] MuI._0017_ MuI._3396_ MuI.a_operand\[17\] vssd1 vssd1
+ vccd1 vccd1 MuI._0742_ sky130_fd_sc_hd__a22oi_2
X_09893_ _02530_ _02544_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__nand2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A1 _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6738_ MuI._2653_ MuI._2654_ vssd1 vssd1 vccd1 vccd1 MuI._2655_ sky130_fd_sc_hd__nor2_1
XFILLER_112_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__B2 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _06544_ _04778_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__nand2_1
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__B1 _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A1_N _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06849__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6669_ MuI._0549_ MuI._2578_ vssd1 vssd1 vccd1 vccd1 MuI._2579_ sky130_fd_sc_hd__xnor2_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ _01391_ _01392_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__nand2_1
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07726_ _03324_ _04316_ _00127_ _00126_ _04380_ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__a32o_1
XFILLER_66_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__B1 _04368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _00273_ _00274_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__nor2_1
XFILLER_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12586__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07588_ _00202_ _00203_ _00188_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__a21o_1
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4994__A1 MuI._0725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _01825_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__and3_1
XFILLER_167_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08076__A2 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _01665_ _01672_ _01874_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__o211ai_4
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ _06460_ _05305_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__nand2_1
XFILLER_182_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09189_ _01806_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__inv_2
XANTENNA__10834__A _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ _03959_ _03961_ _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__a21oi_2
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07846__C _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4886__C MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _03902_ _03903_ _03863_ _03864_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a211o_1
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10591__B1 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10102_ _03293_ _05402_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__and2b_1
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11082_ _03692_ _03693_ _03829_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__and3_1
XFILLER_150_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3721__A2 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ _01331_ _02645_ _02694_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a31o_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12883__A2 _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06759__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3799__A MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A a_operand[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6671__A1 MuI._1836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _04792_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12635__A2 _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3949__D MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _02764_ _03671_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__nand2_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1012_ net122 net7 AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0224_ sky130_fd_sc_hd__mux2_1
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _03433_ _03435_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10728__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _05333_ _05469_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and3_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12646__D _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4020_ MuI._3103_ MuI._3104_ MuI._3118_ vssd1 vssd1 vccd1 vccd1 MuI._3120_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13060__A2 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10797_ _03522_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__xnor2_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ AuI.result\[17\] _02732_ _05392_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._510__A AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ _05191_ _05195_ _05320_ _05321_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__a211o_1
XFILLER_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12662__C _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5971_ MuI._1756_ MuI._1757_ vssd1 vssd1 vccd1 vccd1 MuI._1811_ sky130_fd_sc_hd__nor2_1
XFILLER_126_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output92_A net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__A _02815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11418_ _04188_ _04191_ _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__nand3_1
X_12398_ _05246_ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07756__C _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4922_ MuI._0443_ MuI._0448_ MuI._0450_ MuI._0453_ vssd1 vssd1 vccd1 vccd1 MuI._0657_
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ _00345_ _06613_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__a22o_1
XFILLER_180_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._782_ AuI.pe._132_ AuI.pe._320_ AuI.pe._321_ AuI.pe._322_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._323_ sky130_fd_sc_hd__or4_1
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4853_ MuI._0564_ MuI._0566_ MuI._0579_ vssd1 vssd1 vccd1 vccd1 MuI._0582_ sky130_fd_sc_hd__or3_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3804_ MuI._2888_ MuI._2897_ MuI._2903_ vssd1 vssd1 vccd1 vccd1 MuI._2904_ sky130_fd_sc_hd__or3_1
XFILLER_95_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11575__A _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4784_ MuI._0503_ MuI._0505_ MuI._2055_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0506_
+ sky130_fd_sc_hd__and4bb_1
X_13019_ _05911_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06890_ _04240_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__buf_4
XANTENNA__10334__B1 _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6523_ MuI._2416_ MuI._2409_ MuI._2415_ MuI._2417_ vssd1 vssd1 vccd1 vccd1 MuI._2419_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3735_ MuI._2809_ MuI._2834_ vssd1 vssd1 vccd1 vccd1 MuI._2835_ sky130_fd_sc_hd__or2b_1
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6111__B1 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07491__C _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6454_ MuI._1958_ MuI._1961_ MuI._2342_ vssd1 vssd1 vccd1 vccd1 MuI._2343_ sky130_fd_sc_hd__a21oi_1
XMuI._3666_ MuI._2671_ vssd1 vssd1 vccd1 vccd1 MuI._2682_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._3502__A MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _00902_ _00903_ _00904_ _00874_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__a22oi_2
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5405_ MuI._1187_ MuI._1188_ vssd1 vssd1 vccd1 vccd1 MuI._1189_ sky130_fd_sc_hd__nor2_1
XFILLER_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6385_ MuI._2250_ MuI._2252_ MuI._2266_ vssd1 vssd1 vccd1 vccd1 MuI._2267_ sky130_fd_sc_hd__or3_1
X_07511_ _00123_ _00128_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__xor2_4
XMuI._3597_ MuI._0581_ MuI._0746_ MuI._0801_ MuI._1153_ vssd1 vssd1 vccd1 vccd1 MuI._1923_
+ sky130_fd_sc_hd__and4_1
X_08491_ _00889_ _01106_ _01107_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5336_ MuI._1110_ MuI._1112_ vssd1 vssd1 vccd1 vccd1 MuI._1113_ sky130_fd_sc_hd__or2_1
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4036__C MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._404__B AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ _00058_ _00059_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__nand2_1
XFILLER_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5267_ MuI._0914_ MuI._0916_ MuI._0915_ vssd1 vssd1 vccd1 vccd1 MuI._1037_ sky130_fd_sc_hd__o21bai_1
X_07373_ _06659_ _06660_ _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a21oi_2
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4218_ MuI._1472_ MuI._2843_ MuI._2874_ MuI._2876_ vssd1 vssd1 vccd1 vccd1 MuI._3318_
+ sky130_fd_sc_hd__and4_1
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09112_ _01727_ _01728_ _01719_ _01723_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a211oi_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5198_ MuI._0954_ MuI._0956_ MuI._0960_ vssd1 vssd1 vccd1 vccd1 MuI._0961_ sky130_fd_sc_hd__a21o_1
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4149_ MuI._3244_ MuI._3248_ vssd1 vssd1 vccd1 vccd1 MuI._3249_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ _01646_ _01585_ _01659_ _01660_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__o211ai_2
XFILLER_176_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07666__C _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07385__D _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09945_ _02596_ _02607_ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__or2_1
XANTENNA_AuI.pe._546__A1 AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0908__A AuI._0127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08778__B _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _02118_ _04057_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a21boi_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5611__B MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _01442_ _01443_ _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__o21bai_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _00878_ _00301_ _00259_ _00877_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__a22oi_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__B1 _04631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07709_ _00319_ _00326_ vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__xor2_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _01245_ _01268_ _01263_ _01267_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__o211ai_4
XFILLER_26_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _03439_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__nand2_1
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07203__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09121__C _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _03365_ _03363_ _03364_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__nand3_1
XFILLER_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6169__B1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5058__B MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _03831_ _05842_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
X_10582_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _00237_ _00096_ _05756_ _00785_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__and4_1
XFILLER_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _00502_ _04918_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nand2_2
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3942__A2 MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1630_ AuI._0693_ AuI._0791_ AuI._0795_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0796_
+ sky130_fd_sc_hd__o22a_1
X_11203_ _00727_ _00197_ _00421_ _00728_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a22oi_1
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12183_ _02751_ _04901_ _05002_ _05016_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__a211o_4
XFILLER_135_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5505__C MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1073__A2 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6341__B1 MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1561_ AuI.pe.Significand\[7\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0740_
+ sky130_fd_sc_hd__or2_1
X_11134_ _00345_ _04725_ _03883_ _03885_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__nand4_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0820__A2 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0818__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08509__B1 _00896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11065_ _03810_ _03811_ _03634_ _03638_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o211ai_1
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1492_ AuI._0613_ AuI._0614_ AuI._0620_ AuI._0677_ AuI._0615_ vssd1 vssd1 vccd1
+ vccd1 AuI._0678_ sky130_fd_sc_hd__o221a_1
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09182__B1 _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10016_ _01876_ _01878_ _02684_ _02674_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a211oi_2
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4418__A MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3520_ MuI._1043_ MuI._0471_ MuI._1054_ MuI._1065_ vssd1 vssd1 vccd1 vccd1 MuI._1076_
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12069__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4137__B MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3451_ MuI.a_operand\[24\] MuI.b_operand\[24\] vssd1 vssd1 vccd1 vccd1 MuI._0317_
+ sky130_fd_sc_hd__or2_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10619__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _04781_ _04782_ _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nand3_1
XMuI._6170_ MuI._0328_ MuI._2894_ MuI._2802_ MuI._2803_ vssd1 vssd1 vccd1 vccd1 MuI._2030_
+ sky130_fd_sc_hd__and4_1
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13115__A _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10918_ _03652_ _03478_ _03653_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o21ai_4
XFILLER_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5121_ MuI._0873_ MuI._0874_ MuI._0875_ vssd1 vssd1 vccd1 vccd1 MuI._0876_ sky130_fd_sc_hd__or3_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ _02965_ _04854_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__nand2_1
XFILLER_177_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _00086_ _00462_ _05025_ _06623_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand4_1
XFILLER_158_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5052_ MuI._0168_ MuI._0228_ vssd1 vssd1 vccd1 vccd1 MuI._0800_ sky130_fd_sc_hd__nand2_1
XFILLER_201_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06952__A _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4003_ MuI._3100_ MuI._3101_ MuI._3102_ vssd1 vssd1 vccd1 vccd1 MuI._3103_ sky130_fd_sc_hd__and3_1
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12519_ _03134_ _05360_ _05361_ _05367_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a311o_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11347__A2 _00445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5954_ MuI._1790_ MuI._1792_ vssd1 vssd1 vccd1 vccd1 MuI._1793_ sky130_fd_sc_hd__nor2_1
XFILLER_126_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4905_ MuI._0637_ MuI._0638_ vssd1 vssd1 vccd1 vccd1 MuI._0639_ sky130_fd_sc_hd__xnor2_2
XMuI._5885_ MuI._1667_ MuI._1704_ MuI._1702_ vssd1 vssd1 vccd1 vccd1 MuI._1717_ sky130_fd_sc_hd__a21boi_1
XFILLER_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07991_ _00312_ _00606_ _00603_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__and3_1
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4836_ MuI._2605_ MuI._3306_ MuI._2881_ MuI._2852_ vssd1 vssd1 vccd1 vccd1 MuI._0563_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_141_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._765_ AuI.pe._211_ AuI.pe._002_ AuI.pe._173_ AuI.pe._393_ AuI.pe._308_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._309_ sky130_fd_sc_hd__a221o_1
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5712__A MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _02304_ _02306_ _02305_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a21o_1
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06942_ _04800_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__and3_1
XANTENNA__10307__B1 _00698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4767_ MuI._0288_ MuI._0287_ vssd1 vssd1 vccd1 vccd1 MuI._0487_ sky130_fd_sc_hd__nor2_1
XAuI.pe._696_ AuI.pe._059_ AuI.pe._397_ AuI.pe._213_ AuI.pe._055_ AuI.pe._242_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._243_ sky130_fd_sc_hd__a221o_1
X_09661_ _02294_ _02295_ _02299_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__nand3_1
X_06873_ _04057_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__buf_4
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11455__D _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3718_ MuI._2817_ MuI._2363_ MuI._2812_ MuI._2815_ vssd1 vssd1 vccd1 vccd1 MuI._2818_
+ sky130_fd_sc_hd__o2bb2a_1
XMuI._6506_ MuI._2044_ MuI._2088_ MuI._2033_ vssd1 vssd1 vccd1 vccd1 MuI._2400_ sky130_fd_sc_hd__o21ba_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08612_ _06583_ _04638_ _00033_ _06585_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a22oi_1
XMuI._4698_ MuI._0407_ MuI._0408_ vssd1 vssd1 vccd1 vccd1 MuI._0411_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._5150__C MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _06560_ _03960_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__nand2_1
XFILLER_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6437_ MuI._2322_ MuI._2323_ vssd1 vssd1 vccd1 vccd1 MuI._2324_ sky130_fd_sc_hd__and2b_1
XMuI._3649_ MuI._2484_ vssd1 vssd1 vccd1 vccd1 MuI._2495_ sky130_fd_sc_hd__buf_2
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _01158_ _01160_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__nor2_1
XANTENNA_AuI.pe._700__B2 AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6368_ MuI._2081_ MuI._2080_ MuI._2076_ vssd1 vssd1 vccd1 vccd1 MuI._2248_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1278__B AuI._0477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _01091_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XFILLER_211_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__A _00734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5319_ MuI._3349_ MuI._3262_ MuI._3397_ MuI._2785_ vssd1 vssd1 vccd1 vccd1 MuI._1094_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07023__A _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6299_ MuI._2170_ MuI._2171_ vssd1 vssd1 vccd1 vccd1 MuI._2172_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07425_ _03002_ _00036_ _00031_ _00034_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_168_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A _00567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__A2 _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3621__A1 MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _06543_ _06552_ _06542_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06862__A _03939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4998__A MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11586__A2 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12075__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07287_ _06582_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__nor2_1
XANTENNA__09595__D _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _01547_ _01627_ _01642_ _01643_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__o211a_1
XFILLER_164_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._767__B2 AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12535__A1 _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12535__B2 _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09928_ _02028_ _02587_ _02336_ _02586_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a211o_1
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4885__B1 MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ _02473_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__nand2_1
XFILLER_74_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6626__A1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4637__B1 MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12870_ _05748_ _05752_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__o21a_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12758__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _02669_ _04607_ _02743_ _02944_ _04542_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a32o_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3796__B MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04499_ _04551_ _04552_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__and3_1
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10278__B _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _03419_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__xnor2_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11683_ _04298_ _04363_ _04477_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o211a_2
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13422_ _02817_ _06315_ _06335_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__o21a_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12223__B1 _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10634_ _06429_ _04251_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nand2_1
XANTENNA__06772__A _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ FuI.Integer\[27\] _04627_ _03675_ _05788_ _06265_ vssd1 vssd1 vccd1 vccd1
+ _06266_ sky130_fd_sc_hd__a221o_1
X_10565_ _03272_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__xor2_1
XANTENNA__10294__A _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0992_ AuI._0031_ AuI._0101_ AuI._0194_ vssd1 vssd1 vccd1 vccd1 AuI._0204_ sky130_fd_sc_hd__nand3_1
XFILLER_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09805__A1_N _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ _05075_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
XANTENNA_AuI.pe._758__A1 AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _06191_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10496_ _00077_ _00059_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nand2_1
XFILLER_170_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12235_ _04917_ _04934_ _05072_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10444__D _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4463__A2_N MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1613_ AuI._0701_ AuI._0781_ AuI._0782_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0783_
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ _04870_ _04871_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nor2_1
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5670_ MuI._1001_ MuI._1000_ vssd1 vssd1 vccd1 vccd1 MuI._1480_ sky130_fd_sc_hd__and2b_1
XAuI._1544_ AuI.pe.Significand\[4\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0726_
+ sky130_fd_sc_hd__or2_1
XFILLER_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11117_ _03658_ _04531_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3679__B2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _00262_ _03071_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nand2_1
XMuI._4621_ MuI._0301_ MuI._0325_ vssd1 vssd1 vccd1 vccd1 MuI._0326_ sky130_fd_sc_hd__or2_1
XAuI.pe._550_ AuI.pe._106_ AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 AuI.pe._107_ sky130_fd_sc_hd__nor2_1
XANTENNA__10460__C _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08211__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07108__A _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11048_ _03785_ _03792_ _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nand3_1
XAuI._1475_ AuI._0392_ AuI._0395_ vssd1 vssd1 vccd1 vccd1 AuI._0661_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._4148__A MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._481_ AuI.pe._044_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[2\] sky130_fd_sc_hd__clkbuf_1
Xinput8 a_operand[12] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_6
XANTENNA__07705__A1 _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4552_ MuI._0238_ MuI._0248_ vssd1 vssd1 vccd1 vccd1 MuI._0250_ sky130_fd_sc_hd__nor2_1
XANTENNA__07705__B2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3503_ MuI._0878_ vssd1 vssd1 vccd1 vccd1 MuI._0889_ sky130_fd_sc_hd__buf_2
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06947__A _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A2 _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4483_ MuI._0038_ MuI._0173_ vssd1 vssd1 vccd1 vccd1 MuI._0175_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6222_ MuI.b_operand\[19\] MuI._2811_ MuI._2840_ MuI._2616_ vssd1 vssd1 vccd1
+ vccd1 MuI._2087_ sky130_fd_sc_hd__and4_1
XFILLER_91_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ _03733_ _05520_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__nand2_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3434_ MuI._0086_ MuI._0097_ MuI._0108_ vssd1 vssd1 vccd1 vccd1 MuI._0130_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07469__B1 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10188__B _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6153_ MuI._2008_ MuI._2009_ MuI._2010_ MuI._0570_ MuI._2583_ vssd1 vssd1 vccd1
+ vccd1 MuI._2012_ sky130_fd_sc_hd__o2111a_1
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5104_ MuI._0851_ MuI._0852_ MuI._0857_ vssd1 vssd1 vccd1 vccd1 MuI._0858_ sky130_fd_sc_hd__a21o_1
XFILLER_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08881__B _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6084_ MuI._1931_ MuI._1935_ vssd1 vssd1 vccd1 vccd1 MuI._1936_ sky130_fd_sc_hd__xnor2_1
X_07210_ _06485_ _06509_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__nand3_2
X_08190_ _00481_ _00521_ _00480_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__a21boi_2
XANTENNA__07778__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5035_ MuI._0673_ MuI._0781_ vssd1 vssd1 vccd1 vccd1 MuI._0782_ sky130_fd_sc_hd__nor2_1
XANTENNA__11568__A2 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ _03593_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4611__A MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__D _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _04327_ _06067_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__and2_1
XFILLER_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10354__D _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6305__B1 MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5937_ MuI._0727_ MuI._1724_ MuI._1726_ MuI._1728_ vssd1 vssd1 vccd1 vccd1 MuI._1774_
+ sky130_fd_sc_hd__or4_1
XFILLER_142_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08402__A _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._817_ AuI.pe.significand\[7\] AuI.pe._273_ AuI.pe._070_ AuI.pe._353_ AuI.pe._355_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._356_ sky130_fd_sc_hd__o311a_1
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5868_ MuI._1622_ MuI._1684_ MuI._1696_ MuI._1697_ vssd1 vssd1 vccd1 vccd1 MuI._1698_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07974_ net123 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__buf_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._748_ AuI.pe._276_ AuI.pe._279_ AuI.pe._289_ AuI.pe._292_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[21\] sky130_fd_sc_hd__o31a_1
XMuI._4819_ MuI._0542_ MuI._0543_ vssd1 vssd1 vccd1 vccd1 MuI._0544_ sky130_fd_sc_hd__xor2_1
X_09713_ _02298_ _02297_ _02296_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07018__A net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06925_ _04618_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[10\] sky130_fd_sc_hd__dlymetal6s2s_1
XMuI._5799_ MuI._1608_ MuI._1620_ MuI._1621_ vssd1 vssd1 vccd1 vccd1 MuI._1622_ sky130_fd_sc_hd__nand3_1
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13454__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._679_ AuI.pe._046_ AuI.pe._397_ AuI.pe._225_ AuI.pe._030_ AuI.pe._226_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._227_ sky130_fd_sc_hd__a221o_1
XFILLER_110_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _02274_ _02276_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__and2b_1
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06856_ _03873_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06857__A _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10700__B1 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11482__B _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4208__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09575_ _02120_ _02121_ _02122_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__and3_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06787_ _03131_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[19\] sky130_fd_sc_hd__clkbuf_2
XANTENNA__10379__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__D _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03217_ _03271_ net132 _06430_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__and4_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ _01071_ _01074_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__or2b_1
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._161_ FuI.a_operand\[31\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07408_ _06576_ _06641_ _00024_ _00025_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__a211o_1
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _00832_ _00831_ _00824_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a21o_1
XFILLER_183_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFuI._092_ FuI._052_ FuI._053_ net105 FuI.a_operand\[7\] vssd1 vssd1 vccd1 vccd1 FuI._019_
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07339_ _06637_ _06638_ _06596_ _06616_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__a211o_1
XFILLER_109_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5347__A1 MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5347__B2 MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ _00771_ _00779_ _00778_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__a21o_1
XFILLER_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12508__B2 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _01547_ _01548_ _01562_ _01563_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__and4bb_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _02967_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI._1028__A2 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__A1 _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _04727_ _04729_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__nand2_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11657__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__C _00471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09127__B _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07573__D _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5071__B MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _05808_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__xnor2_1
XAuI._1260_ AuI._0438_ AuI._0333_ vssd1 vssd1 vccd1 vccd1 AuI._0461_ sky130_fd_sc_hd__nand2_1
XFILLER_19_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06767__A _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A2 _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _05648_ _05651_ _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1191_ AuI._0256_ AuI._0393_ AuI._0394_ AuI._0395_ vssd1 vssd1 vccd1 vccd1 AuI._0397_
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13236__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _04606_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__nand2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12784_ _05599_ _05600_ _05661_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a211oi_2
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11735_ _00237_ _00462_ _06489_ _05498_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__and4_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0831__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07598__A _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _04458_ _04459_ _04448_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _06299_ _06301_ _06314_ _06319_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__a211o_4
XFILLER_128_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ _03288_ _03285_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__and2b_2
XFILLER_155_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ _04232_ _04235_ _04233_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12009__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ _06225_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__xor2_1
X_10548_ _00785_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0975_ AuI._0164_ AuI._0169_ AuI._0186_ vssd1 vssd1 vccd1 vccd1 AuI._0187_ sky130_fd_sc_hd__and3_1
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6840_ MuI._2752_ vssd1 vssd1 vccd1 vccd1 MuI.result\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_109_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13267_ _03755_ _05788_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand3_1
X_10479_ _03045_ _03046_ _03048_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o21bai_1
XMuI._3983_ MuI._3071_ MuI._3080_ vssd1 vssd1 vccd1 vccd1 MuI._3083_ sky130_fd_sc_hd__xnor2_1
XMuI._6771_ MuI._2620_ vssd1 vssd1 vccd1 vccd1 MuI._2691_ sky130_fd_sc_hd__clkinv_2
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12218_ _03228_ _03282_ _05509_ _05574_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and4_1
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08222__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _05947_ _06041_ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__or3_1
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5722_ MuI._1534_ MuI._1535_ MuI._1519_ vssd1 vssd1 vccd1 vccd1 MuI._1537_ sky130_fd_sc_hd__a21o_1
XFILLER_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _04977_ _04978_ _04942_ _04808_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__o211a_1
XAuI.pe._602_ AuI.pe._029_ AuI.pe._133_ AuI.pe._150_ AuI.pe._030_ AuI.pe._155_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._156_ sky130_fd_sc_hd__a221o_1
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4322__A_N MuI._3418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5653_ MuI._1062_ MuI._1179_ vssd1 vssd1 vccd1 vccd1 MuI._1462_ sky130_fd_sc_hd__nor2_1
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1527_ AuI._0653_ AuI._0654_ AuI._0656_ vssd1 vssd1 vccd1 vccd1 AuI._0711_ sky130_fd_sc_hd__a21o_1
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5412__D MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._533_ AuI.pe._063_ AuI.pe._042_ AuI.pe._079_ AuI.pe._029_ AuI.pe._091_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._092_ sky130_fd_sc_hd__a221o_1
XMuI._4604_ MuI._0303_ MuI._0307_ vssd1 vssd1 vccd1 vccd1 MuI._0308_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4309__C MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5584_ MuI._3269_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._1386_ sky130_fd_sc_hd__nand2_1
X_06710_ _02302_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__and3_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1458_ AuI._0634_ AuI._0643_ vssd1 vssd1 vccd1 vccd1 AuI._0644_ sky130_fd_sc_hd__or2b_1
X_07690_ _00305_ _00307_ vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__and2b_1
XFILLER_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4535_ MuI._0230_ MuI._0231_ vssd1 vssd1 vccd1 vccd1 MuI._0232_ sky130_fd_sc_hd__nor2_1
XAuI.pe._464_ AuI.pe._028_ vssd1 vssd1 vccd1 vccd1 AuI.pe._029_ sky130_fd_sc_hd__buf_2
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3718__A1_N MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10199__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1389_ AuI._0578_ AuI._0579_ vssd1 vssd1 vccd1 vccd1 AuI._0580_ sky130_fd_sc_hd__nand2_2
XANTENNA_MuI._4606__A MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4466_ MuI._2066_ MuI._2895_ vssd1 vssd1 vccd1 vccd1 MuI._0156_ sky130_fd_sc_hd__nand2_1
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09360_ _01971_ _01976_ _01972_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nand3_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6205_ MuI._0592_ MuI._2860_ MuI._2068_ vssd1 vssd1 vccd1 vccd1 MuI._2069_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08311_ _00928_ _00608_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__xnor2_2
XMuI._4397_ MuI._2704_ MuI._2649_ MuI._2495_ MuI._2773_ vssd1 vssd1 vccd1 vccd1 MuI._0080_
+ sky130_fd_sc_hd__and4_1
XFILLER_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _01908_ _01804_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6136_ MuI._1917_ MuI._1992_ vssd1 vssd1 vccd1 vccd1 MuI._1993_ sky130_fd_sc_hd__xnor2_2
XFILLER_178_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10188__A_N _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _00555_ _00566_ _00565_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__a21boi_2
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10461__A2 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10646__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6067_ MuI._1843_ MuI._1845_ MuI._1916_ vssd1 vssd1 vccd1 vccd1 MuI._1917_ sky130_fd_sc_hd__o21ai_2
XFILLER_193_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07301__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__D _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _06463_ net111 net28 net29 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._4341__A MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5018_ MuI._0760_ MuI._0761_ MuI._0707_ MuI._0762_ vssd1 vssd1 vccd1 vccd1 MuI._0763_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout124_A net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07124_ _05992_ _06056_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__and2_1
XANTENNA__07614__B1 _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07055_ net3 vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__buf_2
XANTENNA__11758__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5172__A MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10812__D _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4304__A2 MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _00571_ _00574_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__or2b_1
XANTENNA__13466__A2 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11493__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06908_ _04434_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__buf_4
XANTENNA__07690__B _00307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11477__A1 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07888_ net112 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__buf_2
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _02258_ _02263_ _02214_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a211o_1
XFILLER_71_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06839_ _03680_ _03690_ _03185_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__and3_1
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _02104_ _02101_ _02103_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a21o_1
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ _00892_ _00893_ _00896_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__o21a_1
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _02113_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nor2_1
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _04300_ _04301_ _04142_ _04145_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a211oi_4
XFILLER_200_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._144_ FuI._006_ net150 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[15\] sky130_fd_sc_hd__dlxtn_1
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _04034_ _04037_ _04036_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__o21bai_1
XFILLER_184_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._075_ FuI._041_ vssd1 vssd1 vccd1 vccd1 FuI._014_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10275__C _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _03068_ _03098_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__xnor2_2
XANTENNA_MuI._5066__B MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11382_ _04023_ _04008_ _04153_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__and3_1
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__A2 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ _03669_ _05660_ _05956_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a31o_1
X_10333_ _03023_ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input54_A b_operand[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _05870_ _05873_ _05946_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__or3_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10264_ _00815_ _02703_ _00814_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a21o_1
XFILLER_133_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5082__A MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12901__A1 _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__xor2_1
XANTENNA__12901__B2 _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _04929_ _02916_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__or2b_1
XFILLER_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13094__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1312_ AuI._0494_ AuI._0495_ AuI._0478_ vssd1 vssd1 vccd1 vccd1 AuI._0510_ sky130_fd_sc_hd__or3b_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6048__A2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ _05790_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__xnor2_1
XAuI._1243_ AuI._0437_ AuI._0441_ AuI._0443_ AuI._0444_ vssd1 vssd1 vccd1 vccd1 AuI._0446_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08752__A2_N _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4320_ MuI._3257_ MuI._3419_ vssd1 vssd1 vccd1 vccd1 MuI._3420_ sky130_fd_sc_hd__xor2_2
XANTENNA_MuI._4426__A MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1174_ AuI._0379_ AuI._0380_ vssd1 vssd1 vccd1 vccd1 AuI._0381_ sky130_fd_sc_hd__nand2_2
X_12836_ _05716_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__nor2_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4251_ MuI._2517_ MuI._2786_ MuI._2352_ MuI._2550_ vssd1 vssd1 vccd1 vccd1 MuI._3351_
+ sky130_fd_sc_hd__a22oi_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12968__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08097__B1 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11850__B _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ net61 _05262_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__nand2_1
XANTENNA__10979__B1 _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08636__A2 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4182_ MuI._3255_ MuI._3280_ MuI._3281_ vssd1 vssd1 vccd1 vccd1 MuI._3282_ sky130_fd_sc_hd__a21oi_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11718_ _00058_ _03071_ _04514_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a22o_1
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10443__A2 _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ _05567_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nand2_1
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput11 a_operand[15] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_6
XFILLER_128_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11649_ _04261_ _04263_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a21oi_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 a_operand[25] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_4
Xinput33 a_operand[6] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_6
Xinput44 b_operand[16] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_8
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput55 b_operand[26] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_6
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6787__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput66 b_operand[7] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_6
XFILLER_183_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13319_ _06108_ _06228_ _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__o21a_1
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10482__A _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0958_ net119 net13 AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0170_ sky130_fd_sc_hd__mux2_1
XMuI._6823_ MuI._2742_ vssd1 vssd1 vccd1 vccd1 MuI.result\[3\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_MuI._4534__A2 MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__B1 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0889_ AuI._0108_ net55 net131 AuI._0107_ vssd1 vssd1 vccd1 vccd1 AuI._0109_
+ sky130_fd_sc_hd__a2bb2o_1
XMuI._6754_ MuI._2656_ MuI._2661_ MuI._2665_ vssd1 vssd1 vccd1 vccd1 MuI._2673_ sky130_fd_sc_hd__a21oi_1
XMuI._3966_ MuI._0581_ MuI._2898_ MuI._3058_ MuI._3065_ vssd1 vssd1 vccd1 vccd1 MuI._3066_
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _01474_ _01477_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__xnor2_2
XFILLER_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5705_ MuI._1036_ MuI._1045_ MuI._1044_ vssd1 vssd1 vccd1 vccd1 MuI._1519_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._6287__A2 MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _00419_ _00420_ _00427_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4298__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3897_ MuI._2983_ MuI._2985_ MuI._2984_ vssd1 vssd1 vccd1 vccd1 MuI._2997_ sky130_fd_sc_hd__o21bai_1
XMuI._6685_ MuI._2596_ vssd1 vssd1 vccd1 vccd1 MuI._2597_ sky130_fd_sc_hd__inv_2
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08791_ _03174_ _03895_ _01405_ _01406_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5636_ MuI._1438_ MuI._1442_ vssd1 vssd1 vccd1 vccd1 MuI._1443_ sky130_fd_sc_hd__and2_1
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07742_ _00341_ _00333_ _00359_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__o21a_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._516_ AuI.pe._385_ AuI.pe._386_ vssd1 vssd1 vccd1 vccd1 AuI.pe._076_ sky130_fd_sc_hd__nor2_1
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5567_ MuI._1364_ MuI._1359_ MuI._1341_ MuI._1366_ vssd1 vssd1 vccd1 vccd1 MuI._1367_
+ sky130_fd_sc_hd__o211a_1
X_07673_ _00289_ _06433_ _04176_ _00290_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a22oi_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._447_ AuI.pe.significand\[0\] vssd1 vssd1 vccd1 vccd1 AuI.pe._014_ sky130_fd_sc_hd__buf_2
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4518_ MuI._0210_ MuI._0211_ MuI._0212_ vssd1 vssd1 vccd1 vccd1 MuI._0213_ sky130_fd_sc_hd__o21ba_1
X_09412_ _02021_ _02028_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a211oi_2
XANTENNA_AuI._0923__A1 net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5498_ MuI._1233_ MuI._1286_ MuI._1282_ MuI._1284_ vssd1 vssd1 vccd1 vccd1 MuI._1291_
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12408__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10682__A2 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3597__D MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4449_ MuI._0128_ MuI._0129_ vssd1 vssd1 vccd1 vccd1 MuI._0137_ sky130_fd_sc_hd__and2b_1
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09343_ _01959_ _01960_ _01844_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a21o_1
XANTENNA__12959__B2 _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08772__D _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _01890_ _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__xor2_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6119_ MuI._1972_ MuI._1973_ vssd1 vssd1 vccd1 vccd1 MuI._1974_ sky130_fd_sc_hd__nor2_2
XFILLER_21_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07031__A _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08225_ _00840_ _00841_ _00842_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__o21ba_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08156_ _06565_ _06516_ _05563_ _05638_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__nand4_1
XFILLER_181_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07107_ _06417_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[22\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ _00491_ _00493_ _00703_ _00704_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__a211oi_1
XFILLER_164_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _05831_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__clkbuf_4
XFILLER_162_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._140__146 vssd1 vssd1 vccd1 vccd1 FuI._140__146/HI net146 sky130_fd_sc_hd__conb_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11147__B1 _03879_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08989_ _01345_ _01346_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__xor2_1
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ _02760_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4246__A MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11870__A1 _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ _03612_ _03613_ _03605_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a21o_1
XFILLER_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _02852_ _05382_ _05379_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a21o_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or2b_1
XFILLER_185_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _04121_ _04126_ _04283_ _04284_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a211o_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12483_ _05228_ _05230_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a211o_2
XFILLER_138_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFuI._127_ net105 FuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 FuI._032_ sky130_fd_sc_hd__and2_1
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _00088_ _06568_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__nand2_4
XANTENNA__06780__A _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0812_ net51 net19 vssd1 vssd1 vccd1 vccd1 AuI._0032_ sky130_fd_sc_hd__xor2_1
XFILLER_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _04134_ _04135_ _03983_ _03985_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__a211o_1
XFILLER_125_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13104_ _03346_ _05467_ _02744_ _04627_ FuI.Integer\[23\] vssd1 vssd1 vccd1 vccd1
+ _06006_ sky130_fd_sc_hd__a32o_1
XANTENNA_MuI._4516__A2 MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10316_ _00716_ _00717_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__nand2_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ _04059_ _04060_ _04055_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__a21o_1
XMuI._3820_ MuI._2704_ MuI._2627_ MuI._2919_ MuI._2916_ vssd1 vssd1 vccd1 vccd1 MuI._2920_
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08203__C _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13035_ _03293_ _05402_ _02742_ _02943_ _05338_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a32o_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ MuI.result\[1\] _02739_ _02719_ _04068_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__a221o_1
XFILLER_121_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12886__B1 _05754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3751_ MuI._2850_ vssd1 vssd1 vccd1 vccd1 MuI._2851_ sky130_fd_sc_hd__buf_4
XFILLER_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11845__B _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _04607_ _02669_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__or2b_1
XFILLER_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6470_ MuI._2351_ MuI._2359_ vssd1 vssd1 vccd1 vccd1 MuI._2360_ sky130_fd_sc_hd__xnor2_1
XMuI._3682_ MuI._2572_ MuI._2743_ MuI._2736_ vssd1 vssd1 vccd1 vccd1 MuI._2782_ sky130_fd_sc_hd__a21o_1
XFILLER_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13118__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09315__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5421_ MuI._1203_ MuI._1205_ vssd1 vssd1 vccd1 vccd1 MuI._1206_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07116__A _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5352_ MuI._1095_ MuI._1094_ MuI._1093_ vssd1 vssd1 vccd1 vccd1 MuI._1130_ sky130_fd_sc_hd__o21ai_1
XAuI._1226_ AuI._0396_ AuI._0416_ vssd1 vssd1 vccd1 vccd1 AuI._0430_ sky130_fd_sc_hd__nor2_1
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4303_ MuI._3402_ vssd1 vssd1 vccd1 vccd1 MuI._3403_ sky130_fd_sc_hd__buf_2
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5283_ MuI._1014_ MuI._1015_ MuI._1052_ MuI._1053_ vssd1 vssd1 vccd1 vccd1 MuI._1055_
+ sky130_fd_sc_hd__or4_1
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1157_ AuI._0328_ AuI._0326_ AuI._0347_ AuI._0348_ vssd1 vssd1 vccd1 vccd1 AuI._0365_
+ sky130_fd_sc_hd__o31a_2
X_12819_ _00278_ _00279_ _06537_ _05756_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__and4_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4234_ MuI._3218_ MuI._3217_ vssd1 vssd1 vccd1 vccd1 MuI._3334_ sky130_fd_sc_hd__nor2_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1088_ net16 net48 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0299_ sky130_fd_sc_hd__mux2_1
XFILLER_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09282__A2 _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4165_ MuI._3264_ MuI._2883_ MuI._3186_ vssd1 vssd1 vccd1 vccd1 MuI._3265_ sky130_fd_sc_hd__a21o_1
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ _00625_ _00626_ _00627_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__o21bai_1
XMuI._4096_ MuI._3188_ MuI._3194_ MuI._3195_ vssd1 vssd1 vccd1 vccd1 MuI._3196_ sky130_fd_sc_hd__a21bo_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09034__A2 _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06690__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08793__A1 _01407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _02592_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__clkinv_2
XFILLER_171_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3715__B1 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6806_ MuI._2678_ MuI._2727_ MuI._2728_ MuI._2729_ vssd1 vssd1 vccd1 vccd1 MuI._2730_
+ sky130_fd_sc_hd__and4_1
XFILLER_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08912_ _01510_ _01511_ _01528_ _01529_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o211ai_2
XFILLER_98_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4998_ MuI._2605_ MuI.b_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._0741_ sky130_fd_sc_hd__nand2_1
X_09892_ _02522_ _02523_ _02549_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a21o_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6737_ MuI._2645_ MuI._2650_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2654_ sky130_fd_sc_hd__mux2_1
XFILLER_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A2 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3949_ MuI._1461_ MuI._2055_ MuI._2693_ MuI._2638_ vssd1 vssd1 vccd1 vccd1 MuI._3049_
+ sky130_fd_sc_hd__and4_1
X_08843_ _01455_ _01456_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a21o_1
XFILLER_100_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__B2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6668_ MuI._0550_ MuI._2573_ MuI._0547_ vssd1 vssd1 vccd1 vccd1 MuI._2578_ sky130_fd_sc_hd__a21oi_1
XFILLER_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ _01382_ _01387_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12629__B1 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5619_ MuI._1391_ MuI._1390_ vssd1 vssd1 vccd1 vccd1 MuI._1424_ sky130_fd_sc_hd__or2b_1
XANTENNA__07026__A _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _00319_ _00326_ _00342_ vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a21oi_2
XMuI._6599_ MuI._0174_ MuI._2500_ MuI._2501_ vssd1 vssd1 vccd1 vccd1 MuI._2502_ sky130_fd_sc_hd__a21o_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07656_ _03335_ _04186_ _00268_ _00269_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06865__A _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07587_ _00007_ _00016_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__nand2_1
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10387__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _01825_ _01827_ _01826_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a21oi_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _01866_ _01867_ _01873_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__or3_2
XFILLER_194_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12806__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13357__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ _00627_ _00626_ _00625_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _01801_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__and2b_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10834__B _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08139_ _06578_ _06579_ _05370_ _05434_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__and4_1
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07846__D _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11150_ _03863_ _03864_ _03902_ _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__o211ai_4
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4886__D MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0832__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ _02757_ _02760_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__nand3_1
XANTENNA__10850__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _03692_ _03693_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10032_ _02695_ _02696_ _02699_ _01331_ _02701_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a221o_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12883__A3 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3799__B MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6175__B MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A a_operand[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11983_ _04799_ _04801_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nor2_1
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _02764_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__or2_1
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06775__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1011_ AuI._0143_ AuI._0204_ vssd1 vssd1 vccd1 vccd1 AuI._0223_ sky130_fd_sc_hd__nand2_2
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _03439_ _03440_ _03463_ _03464_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__and4_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10297__A _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _05466_ _05468_ _05421_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _02965_ _04380_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nand2_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ _05134_ _03675_ _04642_ _04994_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a221o_1
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12466_ _05309_ _05171_ _05319_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__nor3_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5970_ MuI._1768_ MuI._1794_ vssd1 vssd1 vccd1 vccd1 MuI._1810_ sky130_fd_sc_hd__or2_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _03013_ _05456_ _04189_ _04190_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__nand4_1
XANTENNA__12662__D _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13120__B _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12397_ _02398_ _02584_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nor2_1
XANTENNA__12017__A _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07756__D net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4921_ MuI._0654_ MuI._0655_ vssd1 vssd1 vccd1 vccd1 MuI._0656_ sky130_fd_sc_hd__xor2_2
XFILLER_141_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output85_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ _03389_ _02984_ _00445_ _00550_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nand4_1
XFILLER_180_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._781_ AuI.pe.significand\[5\] AuI.pe.significand\[4\] AuI.pe._388_ AuI.pe._009_
+ AuI.pe._010_ vssd1 vssd1 vccd1 vccd1 AuI.pe._322_ sky130_fd_sc_hd__o2111a_1
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4852_ MuI._0564_ MuI._0566_ MuI._0579_ vssd1 vssd1 vccd1 vccd1 MuI._0580_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11856__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11279_ _04033_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nand3_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3803_ MuI._2899_ MuI._2902_ vssd1 vssd1 vccd1 vccd1 MuI._2903_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13018_ _03831_ _05402_ _05817_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a31o_1
XMuI._4783_ MuI.a_operand\[18\] MuI._0017_ MuI._0018_ MuI.a_operand\[19\] vssd1 vssd1
+ vccd1 vccd1 MuI._0505_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11575__B _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__A1 _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10334__B2 _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6522_ MuI._2264_ MuI._2399_ MuI._2414_ vssd1 vssd1 vccd1 vccd1 MuI._2417_ sky130_fd_sc_hd__o21bai_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6111__A1 MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3734_ MuI._2809_ MuI._2810_ MuI._2833_ vssd1 vssd1 vccd1 vccd1 MuI._2834_ sky130_fd_sc_hd__or3_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6111__B2 MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07491__D _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6453_ MuI._1957_ MuI._1926_ vssd1 vssd1 vccd1 vccd1 MuI._2342_ sky130_fd_sc_hd__and2b_1
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3665_ MuI._2660_ vssd1 vssd1 vccd1 vccd1 MuI._2671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5404_ MuI._3185_ MuI._2829_ MuI._3246_ MuI._2892_ vssd1 vssd1 vccd1 vccd1 MuI._1188_
+ sky130_fd_sc_hd__a22oi_1
X_07510_ _04369_ _00126_ _00127_ vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__a21bo_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6384_ MuI._2263_ MuI._2265_ vssd1 vssd1 vccd1 vccd1 MuI._2266_ sky130_fd_sc_hd__nand2_1
XMuI._3596_ MuI._1901_ MuI._1890_ vssd1 vssd1 vccd1 vccd1 MuI._1912_ sky130_fd_sc_hd__xor2_1
XFILLER_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08490_ _00889_ _01106_ _01107_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__and3_1
XMuI._5335_ MuI._1107_ MuI._1111_ vssd1 vssd1 vccd1 vccd1 MuI._1112_ sky130_fd_sc_hd__or2_1
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4036__D MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07441_ _00048_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__buf_6
XAuI._1209_ AuI._0344_ AuI._0413_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0414_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13036__B1 _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5266_ MuI._1034_ MuI._1035_ vssd1 vssd1 vccd1 vccd1 MuI._1036_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07372_ _06661_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__xor2_1
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__B1 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4217_ MuI._2066_ MuI._2874_ MuI._2876_ MuI._1483_ vssd1 vssd1 vccd1 vccd1 MuI._3317_
+ sky130_fd_sc_hd__a22oi_1
X_09111_ _01719_ _01723_ _01727_ _01728_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__o211a_1
XMuI._5197_ MuI._0957_ MuI._0958_ MuI._0959_ vssd1 vssd1 vccd1 vccd1 MuI._0960_ sky130_fd_sc_hd__o21bai_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4148_ MuI._3247_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._3248_ sky130_fd_sc_hd__nand2_1
XFILLER_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ _01658_ _01657_ _01562_ _01560_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13311__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4079_ MuI._3176_ MuI._3177_ MuI._3178_ vssd1 vssd1 vccd1 vccd1 MuI._3179_ sky130_fd_sc_hd__o21ba_1
XANTENNA_AuI._1067__A0 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07666__D _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09944_ _02597_ _02606_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09715__B1 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _02216_ _06437_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__nand2_1
XANTENNA_input9_A a_operand[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08140__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__C _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5180__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08826_ _02096_ _02194_ net13 net14 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__and4_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08757_ _06606_ _06601_ _04240_ _00074_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__and4_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _00320_ _00325_ vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__xnor2_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08688_ _01269_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _00095_ _00096_ _04358_ _04434_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__and4_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ _03363_ _03364_ _03365_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__a21o_1
XFILLER_198_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09452__A1_N _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09121__D _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6169__A1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _01885_ _01887_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__nor2_1
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6169__B2 MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ _02952_ _03117_ _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5058__C MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12320_ _00081_ _05756_ _00783_ _03056_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a22oi_1
XFILLER_194_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._146__152 vssd1 vssd1 vccd1 vccd1 FuI._146__152/HI net152 sky130_fd_sc_hd__conb_1
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _05087_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__xnor2_4
XFILLER_170_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__B2 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11202_ _03956_ _03957_ _03958_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__a21o_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _05004_ _05006_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a21o_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1073__A3 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6341__A1 MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _03486_ _04725_ _03883_ _03885_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._6341__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1560_ AuI._0701_ AuI._0733_ AuI._0738_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0739_
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11064_ _03634_ _03638_ _03810_ _03811_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__a211o_1
XAuI._1491_ AuI._0673_ AuI._0675_ AuI._0676_ vssd1 vssd1 vccd1 vccd1 AuI._0677_ sky130_fd_sc_hd__a21o_1
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09182__A1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09182__B2 _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _02671_ _02673_ _02672_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o21a_1
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0834__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3450_ MuI._0262_ MuI._0284_ MuI._0295_ vssd1 vssd1 vccd1 vccd1 MuI._0306_ sky130_fd_sc_hd__a21bo_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4137__C MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10619__A2 _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11966_ _04670_ _04669_ _04668_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21bo_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10917_ _03475_ _03477_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__or2_1
XANTENNA__13115__B _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11897_ _00197_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a21bo_1
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5120_ MuI._0327_ MuI._3402_ MuI._3396_ MuI._2429_ vssd1 vssd1 vccd1 vccd1 MuI._0875_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__B _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848_ _00096_ _05025_ _06623_ _00095_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a22o_1
XMuI._5051_ MuI._0796_ MuI._0798_ vssd1 vssd1 vccd1 vccd1 MuI._0799_ sky130_fd_sc_hd__nor2_1
XFILLER_158_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4002_ MuI._2996_ MuI._3005_ MuI._3004_ vssd1 vssd1 vccd1 vccd1 MuI._3102_ sky130_fd_sc_hd__a21bo_1
X_10779_ _02764_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _04159_ _05369_ _05371_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o31ai_4
XANTENNA_AuI._1384__B AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5265__A MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ _05291_ _05211_ _05300_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4600__C MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4591__B1 MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5953_ MuI._1788_ MuI._1789_ MuI._1771_ MuI._1772_ vssd1 vssd1 vccd1 vccd1 MuI._1792_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4904_ MuI._2817_ MuI._0245_ vssd1 vssd1 vccd1 vccd1 MuI._0638_ sky130_fd_sc_hd__nand2_1
XFILLER_153_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5884_ MuI._1651_ MuI._1664_ MuI._1715_ vssd1 vssd1 vccd1 vccd1 MuI._1716_ sky130_fd_sc_hd__a21o_1
XFILLER_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07990_ _03389_ _03454_ _03873_ _03971_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__and4_1
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4343__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._764_ AuI.pe.significand\[20\] AuI.pe._041_ AuI.pe._305_ AuI.pe._306_ AuI.pe._307_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._308_ sky130_fd_sc_hd__a2111o_1
XMuI._4835_ MuI._2671_ MuI._2895_ vssd1 vssd1 vccd1 vccd1 MuI._0562_ sky130_fd_sc_hd__nand2_1
X_06941_ _04789_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._5712__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._695_ AuI.pe._014_ AuI.pe._012_ vssd1 vssd1 vccd1 vccd1 AuI.pe._242_ sky130_fd_sc_hd__and2_1
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4766_ MuI._0484_ MuI._0481_ vssd1 vssd1 vccd1 vccd1 MuI._0486_ sky130_fd_sc_hd__xnor2_1
X_09660_ _02294_ _02295_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a21o_1
X_06872_ _04046_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__buf_6
XMuI._6505_ MuI._2231_ MuI._2253_ vssd1 vssd1 vccd1 vccd1 MuI._2399_ sky130_fd_sc_hd__nor2_1
XFILLER_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3717_ MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 MuI._2817_ sky130_fd_sc_hd__buf_2
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0840__A_N net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _06578_ _06579_ _00030_ _04703_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__and4_1
XFILLER_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4697_ MuI._0371_ MuI._0373_ vssd1 vssd1 vccd1 vccd1 MuI._0410_ sky130_fd_sc_hd__xor2_1
X_09591_ _02222_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__nand2_1
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5150__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6436_ MuI._2313_ MuI._2315_ MuI._2321_ vssd1 vssd1 vccd1 vccd1 MuI._2323_ sky130_fd_sc_hd__or3b_1
XMuI._3648_ MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 MuI._2484_ sky130_fd_sc_hd__clkbuf_4
X_08542_ _01158_ _01159_ _03163_ _06443_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__and4bb_1
XFILLER_211_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6367_ MuI._2081_ MuI._2076_ MuI._2080_ vssd1 vssd1 vccd1 vccd1 MuI._2247_ sky130_fd_sc_hd__and3_1
XANTENNA__07304__A _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3579_ MuI._0724_ MuI._0977_ vssd1 vssd1 vccd1 vccd1 MuI._1725_ sky130_fd_sc_hd__nand2_1
XFILLER_51_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08473_ _01077_ _01078_ _01090_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__and3_1
XFILLER_211_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5318_ MuI._0088_ MuI._3268_ vssd1 vssd1 vccd1 vccd1 MuI._1093_ sky130_fd_sc_hd__nand2_1
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08119__B _00735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _00038_ _00041_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__nor2_1
XFILLER_211_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6298_ MuI._0801_ MuI._1164_ MuI._1043_ MuI._0746_ vssd1 vssd1 vccd1 vccd1 MuI._2171_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_51_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5249_ MuI._0907_ MuI._0910_ MuI._0908_ vssd1 vssd1 vccd1 vccd1 MuI._1017_ sky130_fd_sc_hd__o21bai_1
XFILLER_149_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__A2 _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _06649_ _06650_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._3621__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10243__B1 _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ _06582_ _06586_ _02712_ _04907_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__and4bb_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _01631_ _01632_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__or4bb_1
XFILLER_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07974__A net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12535__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _02586_ _02336_ _02587_ _02028_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__o211ai_4
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4885__A1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13496__B1 _02739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4885__B2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__B_N _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _02467_ _02472_ _02471_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6626__A2 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08809_ _01424_ _01426_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__or2_2
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _02376_ _02382_ _02383_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__or3_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4637__B2 MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4786__A1_N MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _06045_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__buf_2
XFILLER_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07214__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _04549_ _04550_ _04512_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__o21ai_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10702_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__nor2_1
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _04475_ _04476_ _04291_ _04293_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o211ai_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _05788_ _03626_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__or2b_1
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12223__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10633_ _03345_ _03347_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12223__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ MuI.result\[27\] _02737_ _04011_ _02830_ _06263_ vssd1 vssd1 vccd1 vccd1
+ _06265_ sky130_fd_sc_hd__a221o_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _03068_ _03098_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0991_ AuI._0189_ AuI._0192_ AuI._0198_ AuI._0202_ vssd1 vssd1 vccd1 vccd1 AuI._0203_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10785__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _05038_ _05074_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__nor2_1
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13283_ _06128_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__or2_1
X_10495_ _03198_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nor2_1
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12234_ _04915_ _04916_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__or2_1
XANTENNA__07884__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11734__B1 _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1612_ AuI._0769_ AuI._0776_ vssd1 vssd1 vccd1 vccd1 AuI._0782_ sky130_fd_sc_hd__nand2_1
X_12165_ _04996_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__or2_1
XFILLER_111_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11116_ _00059_ _03865_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__a21bo_1
XAuI._1543_ AuI._0701_ AuI._0718_ AuI._0724_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0725_
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12096_ _04921_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__xnor2_1
XMuI._4620_ MuI._0301_ MuI._0302_ MuI._0324_ vssd1 vssd1 vccd1 vccd1 MuI._0325_ sky130_fd_sc_hd__nor3_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08211__C net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10460__D _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _03789_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5251__C MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1474_ AuI._0650_ AuI._0658_ AuI._0659_ AuI._0648_ vssd1 vssd1 vccd1 vccd1 AuI._0660_
+ sky130_fd_sc_hd__and4_1
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4148__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._480_ AuI.pe._034_ AuI.pe._043_ vssd1 vssd1 vccd1 vccd1 AuI.pe._044_ sky130_fd_sc_hd__or2_1
XANTENNA__08902__A1 _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__A2 _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4551_ MuI._0238_ MuI._0248_ vssd1 vssd1 vccd1 vccd1 MuI._0249_ sky130_fd_sc_hd__and2_1
Xinput9 a_operand[13] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_4
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13239__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3502_ MuI._0867_ vssd1 vssd1 vccd1 vccd1 MuI._0878_ sky130_fd_sc_hd__buf_2
XMuI._4482_ MuI._0040_ MuI._0039_ vssd1 vssd1 vccd1 vccd1 MuI._0173_ sky130_fd_sc_hd__nor2_1
XFILLER_92_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6221_ MuI._2053_ MuI._2085_ vssd1 vssd1 vccd1 vccd1 MuI._2086_ sky130_fd_sc_hd__nor2_1
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12998_ _05889_ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__xor2_1
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3433_ MuI._0086_ MuI._0097_ MuI._0108_ vssd1 vssd1 vccd1 vccd1 MuI._0119_ sky130_fd_sc_hd__and3_1
XANTENNA__07124__A _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07469__A1 _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07469__B2 _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4164__A MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _03315_ _04641_ _04651_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a211o_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6152_ MuI._0482_ MuI._0493_ MuI._2006_ vssd1 vssd1 vccd1 vccd1 MuI._2010_ sky130_fd_sc_hd__a21bo_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06963__A _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5103_ MuI._0853_ MuI._0854_ MuI._0855_ vssd1 vssd1 vccd1 vccd1 MuI._0857_ sky130_fd_sc_hd__o21bai_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6083_ MuI._1932_ MuI._1933_ vssd1 vssd1 vccd1 vccd1 MuI._1935_ sky130_fd_sc_hd__nor2_1
XANTENNA__07778__B _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5034_ MuI._0740_ MuI._0778_ MuI._0780_ vssd1 vssd1 vccd1 vccd1 MuI._0781_ sky130_fd_sc_hd__a21oi_2
XFILLER_186_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07140_ _06438_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__A1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3508__A MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07071_ _06181_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_118_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07794__A _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__B _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6305__A1 MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5936_ MuI._1724_ vssd1 vssd1 vccd1 vccd1 MuI._1773_ sky130_fd_sc_hd__inv_2
XANTENNA_MuI._6305__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._816_ AuI.pe._378_ AuI.pe._354_ AuI.pe._380_ vssd1 vssd1 vccd1 vccd1 AuI.pe._355_
+ sky130_fd_sc_hd__or3b_1
XANTENNA__12205__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__B _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5867_ MuI._1687_ MuI._1688_ MuI._1695_ vssd1 vssd1 vccd1 vccd1 MuI._1697_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _00262_ _04316_ _00257_ _00258_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_MuI._4339__A MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._747_ AuI.pe._290_ AuI.pe._291_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._292_
+ sky130_fd_sc_hd__a21o_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4818_ MuI._0409_ MuI._0410_ vssd1 vssd1 vccd1 vccd1 MuI._0543_ sky130_fd_sc_hd__xnor2_1
X_09712_ _02298_ _02296_ _02297_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__or3_1
X_06924_ _04607_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__and3_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5798_ MuI._1612_ MuI._1613_ MuI._1619_ vssd1 vssd1 vccd1 vccd1 MuI._1621_ sky130_fd_sc_hd__a21o_1
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._678_ AuI.pe._063_ AuI.pe._164_ AuI.pe._213_ AuI.pe._028_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._226_ sky130_fd_sc_hd__a22o_1
XANTENNA_AuI.pe._426__A AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4749_ MuI._2429_ MuI._3189_ MuI._3190_ MuI._2660_ vssd1 vssd1 vccd1 vccd1 MuI._0467_
+ sky130_fd_sc_hd__a22oi_1
X_09643_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__inv_2
X_06855_ net115 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10700__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ _02204_ _02206_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nand3_2
X_06786_ _03110_ _03121_ _02680_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__and3_1
XFILLER_71_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10379__B _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6419_ MuI._2301_ MuI._2303_ vssd1 vssd1 vccd1 vccd1 MuI._2304_ sky130_fd_sc_hd__and2b_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07034__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _01138_ _01139_ _01141_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._4074__A MuI._3160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__A _03974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08456_ _01071_ _01072_ _01073_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__or3_1
XFILLER_169_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06873__A _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._160_ FuI.a_operand\[30\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[30\] sky130_fd_sc_hd__clkbuf_1
X_07407_ _06676_ _06677_ _00023_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__nor3_4
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _00964_ _00969_ _00963_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._091_ FuI.a_operand\[26\] FuI._037_ net104 FuI.a_operand\[23\] vssd1 vssd1 vccd1
+ vccd1 FuI._053_ sky130_fd_sc_hd__and4_1
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07338_ _06596_ _06616_ _06637_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__o211ai_4
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10767__A1 _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5347__A2 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ _06559_ _06567_ _06569_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__and3_1
XFILLER_164_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12508__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _01622_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a21boi_1
XFILLER_191_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _00677_ _00681_ _00679_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11716__B1 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1028__A3 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__A2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11657__C _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08312__B _00929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3530__A1 MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _05716_ _05719_ _05717_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o21ba_1
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__C _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12852_ _05653_ _05734_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__xnor2_1
XAuI._1190_ AuI._0255_ AuI._0393_ AuI._0394_ AuI._0395_ vssd1 vssd1 vccd1 vccd1 AuI._0396_
+ sky130_fd_sc_hd__and4_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3600__B MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _03820_ _04607_ _04443_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a31o_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12783_ _05658_ _05659_ _05555_ _05557_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__o211a_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _03099_ _06666_ _00398_ _03056_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__a22oi_2
XFILLER_70_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06783__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11665_ _04448_ _04458_ _04459_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and3_2
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07871__A1 _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _02817_ _06317_ _06318_ _02750_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__o211a_1
X_10616_ _03328_ _03299_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__and2b_1
XFILLER_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11596_ _04239_ _04237_ _04238_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__and3_1
XFILLER_195_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12009__B _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13335_ _06244_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__xnor2_1
X_10547_ _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and2_1
XFILLER_109_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0974_ net49 net17 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0186_ sky130_fd_sc_hd__mux2_1
XFILLER_155_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _06173_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10478_ _03019_ _03039_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nor2_1
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6770_ MuI._2617_ MuI._2687_ MuI._2689_ vssd1 vssd1 vccd1 vccd1 MuI._2690_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI.pe._600__B2 AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _00727_ _03051_ _03071_ _00728_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a22oi_1
XMuI._3982_ MuI._3028_ MuI._3030_ vssd1 vssd1 vccd1 vccd1 MuI._3082_ sky130_fd_sc_hd__xor2_2
XFILLER_124_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or2_1
XFILLER_97_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5721_ MuI._1519_ MuI._1534_ MuI._1535_ vssd1 vssd1 vccd1 vccd1 MuI._1536_ sky130_fd_sc_hd__nand3_2
XANTENNA__08222__B _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ _04942_ _04808_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a211oi_1
XAuI.pe._601_ AuI.pe._102_ AuI.pe._054_ AuI.pe._151_ AuI.pe._154_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._155_ sky130_fd_sc_hd__a211o_1
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5652_ MuI._1182_ MuI._1236_ MuI._1239_ MuI._1458_ MuI._1459_ vssd1 vssd1 vccd1
+ vccd1 MuI._1460_ sky130_fd_sc_hd__a221oi_4
XAuI._1526_ AuI._0709_ vssd1 vssd1 vccd1 vccd1 AuI._0710_ sky130_fd_sc_hd__buf_2
XFILLER_96_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12079_ _04702_ _04749_ _04858_ _04859_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__a211o_1
XAuI.pe._532_ AuI.pe._056_ AuI.pe._050_ AuI.pe._023_ AuI.pe._072_ AuI.pe._090_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._091_ sky130_fd_sc_hd__a221o_1
XANTENNA__06958__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4603_ MuI._2811_ MuI._3246_ MuI._0305_ MuI._2939_ vssd1 vssd1 vccd1 vccd1 MuI._0307_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5583_ MuI._1353_ MuI._1352_ MuI._1350_ vssd1 vssd1 vccd1 vccd1 MuI._1385_ sky130_fd_sc_hd__o21ai_1
XAuI._1457_ AuI._0462_ AuI._0467_ AuI._0640_ AuI._0642_ vssd1 vssd1 vccd1 vccd1 AuI._0643_
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._463_ AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 AuI.pe._028_ sky130_fd_sc_hd__buf_2
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4534_ MuI._1142_ MuI._0101_ MuI._3246_ MuI._2939_ vssd1 vssd1 vccd1 vccd1 MuI._0231_
+ sky130_fd_sc_hd__a22oi_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1388_ AuI._0258_ AuI._0575_ AuI._0576_ AuI._0577_ vssd1 vssd1 vccd1 vccd1 AuI._0579_
+ sky130_fd_sc_hd__a31o_1
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._667__A1 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4606__B MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4465_ MuI._0151_ MuI._0154_ vssd1 vssd1 vccd1 vccd1 MuI._0155_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6204_ MuI._2008_ MuI._2009_ MuI._2010_ vssd1 vssd1 vccd1 vccd1 MuI._2068_ sky130_fd_sc_hd__o21a_1
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__A1 _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _00609_ _00607_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__or2b_1
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4396_ MuI._2919_ MuI._2495_ MuI._2791_ MuI._2800_ vssd1 vssd1 vccd1 vccd1 MuI._0079_
+ sky130_fd_sc_hd__a22oi_1
X_09290_ _06610_ _03971_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__nand2_1
XFILLER_205_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06693__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6135_ MuI._1990_ MuI._1991_ vssd1 vssd1 vccd1 vccd1 MuI._1992_ sky130_fd_sc_hd__nor2_1
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ _02851_ _04660_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__nand2_1
XFILLER_178_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08935__A2_N _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6066_ MuI._1848_ MuI._1847_ vssd1 vssd1 vccd1 vccd1 MuI._1916_ sky130_fd_sc_hd__or2b_1
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08172_ _02248_ _00153_ _00789_ _02205_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__a22oi_1
XFILLER_193_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09064__B1 _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4341__B MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5017_ MuI._0693_ MuI._0706_ MuI._0700_ MuI._0705_ vssd1 vssd1 vccd1 vccd1 MuI._0762_
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ _06425_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[30\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07614__A1 _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07614__B2 _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5156__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout117_A net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ _06003_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[31\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11758__B _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5919_ MuI._1735_ MuI._1753_ vssd1 vssd1 vccd1 vccd1 MuI._1754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5172__B MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10921__A1 _03509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07956_ _00571_ _00572_ _00573_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__or3_1
XANTENNA__06868__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11493__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06907_ net35 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__buf_4
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07887_ _03722_ _03993_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__nand2_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06838_ _02042_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__clkbuf_2
X_09626_ _02211_ _02213_ _02212_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__o21a_1
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _02104_ _02101_ _02103_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__nand3_1
XFILLER_71_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06769_ net44 vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08508_ _01108_ _01109_ _01111_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__or3_1
X_09488_ _01332_ _02334_ _00082_ _00084_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and4_1
XFILLER_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._450__D_N AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ _01010_ _01012_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__or2b_1
XFILLER_157_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._143_ FuI._005_ net149 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[14\] sky130_fd_sc_hd__dlxtn_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11014__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11450_ _06620_ _03257_ _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a22o_1
XFILLER_177_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._074_ FuI.a_operand\[2\] FuI._040_ vssd1 vssd1 vccd1 vccd1 FuI._041_ sky130_fd_sc_hd__and2_1
X_10401_ _03095_ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10275__D _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ _04023_ _04008_ _04153_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _02815_ _05883_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nor2_1
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ _00077_ _04596_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__nand2_1
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _05870_ _05873_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__o21ai_2
X_10263_ _02935_ _02936_ _02937_ _02947_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__a311o_1
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _02965_ _04854_ _04708_ _04707_ _04983_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a32o_1
XANTENNA__12901__A2 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5082__B MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _02842_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__inv_2
XANTENNA_input47_A b_operand[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5513__D MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1311_ AuI._0507_ AuI._0508_ vssd1 vssd1 vccd1 vccd1 AuI._0509_ sky130_fd_sc_hd__nor2_2
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4707__A MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3611__A MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12904_ _02987_ _05713_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nand2_1
XAuI._1242_ AuI._0437_ AuI._0441_ AuI._0443_ AuI._0444_ vssd1 vssd1 vccd1 vccd1 AuI._0445_
+ sky130_fd_sc_hd__and4_1
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1173_ AuI._0256_ AuI._0377_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0380_ sky130_fd_sc_hd__a21o_1
X_12835_ _00506_ _00676_ _05509_ _05574_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__and4_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0842__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4250_ MuI._3000_ MuI._2754_ MuI._3223_ MuI._3349_ vssd1 vssd1 vccd1 vccd1 MuI._3350_
+ sky130_fd_sc_hd__and4_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08097__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ _05640_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4181_ MuI._3278_ MuI._3279_ vssd1 vssd1 vccd1 vccd1 MuI._3281_ sky130_fd_sc_hd__nor2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _00063_ _00062_ _03425_ _05702_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nand4_1
XFILLER_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11640__A2 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _05348_ _05359_ _05482_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a31o_1
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ _04259_ _04260_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__and2_1
Xinput12 a_operand[16] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput23 a_operand[26] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_6
XFILLER_156_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11928__B1 _04721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 a_operand[7] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
XFILLER_190_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput45 b_operand[17] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_4
X_11579_ _04230_ _04231_ _04236_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nor3b_1
Xinput56 b_operand[27] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_4
Xinput67 b_operand[8] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_4
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _03669_ _05906_ _05981_ _03626_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a22o_1
XAuI._0957_ AuI._0168_ vssd1 vssd1 vccd1 vccd1 AuI._0169_ sky130_fd_sc_hd__clkbuf_2
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10482__B _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6822_ MuI._2713_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2742_ sky130_fd_sc_hd__and2b_1
XFILLER_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _06157_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0888_ AuI._0107_ net131 net23 vssd1 vssd1 vccd1 vccd1 AuI._0108_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11156__B2 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6753_ MuI._2666_ MuI._2670_ vssd1 vssd1 vccd1 vccd1 MuI._2672_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3965_ MuI._3056_ MuI._3057_ vssd1 vssd1 vccd1 vccd1 MuI._3065_ sky130_fd_sc_hd__and2_1
XFILLER_170_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5704_ MuI._1515_ MuI._1517_ vssd1 vssd1 vccd1 vccd1 MuI._1518_ sky130_fd_sc_hd__and2_1
XFILLER_112_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07810_ _00419_ _00420_ _00427_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__nand3_1
XFILLER_85_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6684_ MuI._2591_ MuI._2595_ vssd1 vssd1 vccd1 vccd1 MuI._2596_ sky130_fd_sc_hd__or2_1
XMuI._3896_ MuI._1274_ MuI._2797_ MuI._2931_ MuI._2930_ MuI._2914_ vssd1 vssd1 vccd1
+ vccd1 MuI._2996_ sky130_fd_sc_hd__a32o_1
X_08790_ _03067_ _03110_ _03895_ _03993_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nand4_4
XANTENNA_MuI._4298__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06688__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5635_ MuI._3403_ MuI._0421_ MuI._1414_ MuI._1441_ vssd1 vssd1 vccd1 vccd1 MuI._1442_
+ sky130_fd_sc_hd__and4_1
XAuI._1509_ AuI._0599_ vssd1 vssd1 vccd1 vccd1 AuI._0695_ sky130_fd_sc_hd__buf_2
X_07741_ _00343_ _00358_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__xnor2_2
XAuI.pe._515_ AuI.pe._070_ AuI.pe._073_ AuI.pe._074_ vssd1 vssd1 vccd1 vccd1 AuI.pe._075_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4617__A MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5566_ MuI._1361_ MuI._1363_ MuI._1360_ vssd1 vssd1 vccd1 vccd1 MuI._1366_ sky130_fd_sc_hd__or3_1
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07672_ net113 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__buf_4
XAuI.pe._446_ AuI.pe.significand\[1\] vssd1 vssd1 vccd1 vccd1 AuI.pe._013_ sky130_fd_sc_hd__buf_2
XMuI._4517_ MuI._2799_ MuI._2918_ MuI._2790_ MuI._3223_ vssd1 vssd1 vccd1 vccd1 MuI._0212_
+ sky130_fd_sc_hd__and4_1
X_09411_ _01952_ _01953_ _01954_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__and3_1
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5497_ MuI._1183_ MuI._1235_ MuI._1288_ MuI._1289_ vssd1 vssd1 vccd1 vccd1 MuI._1290_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12408__B2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4448_ MuI._0134_ MuI._0135_ vssd1 vssd1 vccd1 vccd1 MuI._0136_ sky130_fd_sc_hd__xnor2_1
X_09342_ _01765_ _01768_ _01843_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a21o_1
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07312__A _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4379_ MuI._3344_ MuI._3343_ vssd1 vssd1 vccd1 vccd1 MuI._0061_ sky130_fd_sc_hd__nor2_1
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11092__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _02474_ _00089_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__nand2_2
XFILLER_166_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6118_ MuI._0779_ MuI._2802_ MuI._2803_ MuI._2894_ vssd1 vssd1 vccd1 vccd1 MuI._1973_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ _02420_ _06513_ _05025_ _05101_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and4_1
XFILLER_178_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6049_ MuI._1895_ MuI._1896_ vssd1 vssd1 vccd1 vccd1 MuI._1897_ sky130_fd_sc_hd__nor2_1
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _06663_ _00398_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__nand2_1
XFILLER_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11395__B2 _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _05402_ _06414_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__and2_1
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _00701_ _00702_ _00692_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ _05820_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0927__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08988_ _01603_ _01604_ _01602_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a21o_1
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3497__B1 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07939_ _06610_ _04725_ _00038_ _00556_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _03686_ _03687_ _02928_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._5238__A1 MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5238__B2 MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _06488_ _04294_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__and2_1
XFILLER_204_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10881_ _03605_ _03612_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__nand3_1
XFILLER_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__A2 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09421__B _01881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ _02752_ _05384_ _05385_ _05486_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__a31o_2
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08318__A _00934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _05408_ _05409_ _05410_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__a21o_1
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4749__B1 MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11502_ _04281_ _04282_ _04271_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12482_ _05335_ _05336_ _05222_ _05224_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a211oi_2
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._126_ FuI._058_ FuI._026_ FuI._028_ FuI.a_operand\[21\] net105 vssd1 vssd1 vccd1
+ vccd1 FuI._012_ sky130_fd_sc_hd__o2111a_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11433_ _00086_ _00081_ _00412_ _00530_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__and4_1
XFILLER_193_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__B1 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0811_ AuI._0029_ AuI._0030_ vssd1 vssd1 vccd1 vccd1 AuI._0031_ sky130_fd_sc_hd__or2_2
X_11364_ _03983_ _03985_ _04134_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o211ai_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6189__A MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5174__B1 MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13103_ MuI.result\[23\] _02739_ _04642_ _05402_ _06004_ vssd1 vssd1 vccd1 vccd1
+ _06005_ sky130_fd_sc_hd__a221o_1
X_10315_ _00750_ _00764_ _00765_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__nand3_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _04055_ _04059_ _04060_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nand3_1
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13034_ _05402_ _02941_ _02731_ AuI.result\[22\] vssd1 vssd1 vccd1 vccd1 _05931_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10246_ _02216_ _04004_ _02745_ _02931_ FuI.Integer\[1\] vssd1 vssd1 vccd1 vccd1
+ _02932_ sky130_fd_sc_hd__a32o_1
XANTENNA__08203__D _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__B1 _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0837__A net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3750_ MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 MuI._2850_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10177_ _02844_ _02848_ _02853_ _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__or4b_1
XFILLER_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3681_ MuI._2759_ MuI._2780_ vssd1 vssd1 vccd1 vccd1 MuI._2781_ sky130_fd_sc_hd__or2b_1
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13118__B _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__C net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5420_ MuI._1146_ MuI._1204_ vssd1 vssd1 vccd1 vccd1 MuI._1205_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08306__A2 _00922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5351_ MuI._1095_ MuI._1093_ MuI._1094_ vssd1 vssd1 vccd1 vccd1 MuI._1129_ sky130_fd_sc_hd__or3_1
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1225_ AuI._0427_ AuI._0428_ vssd1 vssd1 vccd1 vccd1 AuI._0429_ sky130_fd_sc_hd__xor2_1
XFILLER_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4302_ MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 MuI._3402_ sky130_fd_sc_hd__buf_4
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5282_ MuI._1050_ MuI._1051_ MuI._0924_ MuI._1016_ vssd1 vssd1 vccd1 vccd1 MuI._1053_
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1156_ AuI._0362_ AuI._0363_ vssd1 vssd1 vccd1 vccd1 AuI._0364_ sky130_fd_sc_hd__and2b_2
X_12818_ _03443_ _05702_ _03247_ _00290_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__a22oi_1
XANTENNA__09267__B1 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4233_ MuI._3331_ MuI._3329_ vssd1 vssd1 vccd1 vccd1 MuI._3333_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1087_ AuI._0252_ AuI._0297_ vssd1 vssd1 vccd1 vccd1 AuI._0298_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12810__A1 _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ _05613_ _05622_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__and3_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4164_ MuI._0570_ MuI._2886_ vssd1 vssd1 vccd1 vccd1 MuI._3264_ sky130_fd_sc_hd__nand2_1
XFILLER_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06971__A _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11589__A _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4095_ MuI._2878_ MuI._3187_ MuI._3183_ vssd1 vssd1 vccd1 vccd1 MuI._3195_ sky130_fd_sc_hd__nand3_1
XFILLER_129_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08242__A1 _00555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3516__A MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08793__A2 _01409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09960_ _02617_ _02618_ _02613_ _02623_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a31oi_1
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0841__A1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3715__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6805_ MuI._2656_ MuI._2661_ vssd1 vssd1 vccd1 vccd1 MuI._2729_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3715__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ _01512_ _01513_ _01527_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__nand3_1
XMuI._4997_ MuI._0709_ MuI._0737_ MuI._0739_ vssd1 vssd1 vccd1 vccd1 MuI._0740_ sky130_fd_sc_hd__a21oi_4
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09891_ _02546_ _02548_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__and2b_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6736_ MuI._2650_ MuI._2652_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2653_ sky130_fd_sc_hd__mux2_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3948_ MuI._2916_ MuI._2796_ vssd1 vssd1 vccd1 vccd1 MuI._3048_ sky130_fd_sc_hd__nand2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _01457_ _01458_ _01459_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a21bo_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10196__B_N _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11755__C _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A2 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6667_ MuI._2576_ vssd1 vssd1 vccd1 vccd1 MuI._2577_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3879_ MuI._2974_ MuI._2977_ MuI._2973_ vssd1 vssd1 vccd1 vccd1 MuI._2979_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12629__A1 _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08773_ _03024_ _03982_ _01389_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__a31o_2
XFILLER_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12629__B2 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5618_ MuI._1380_ MuI._1421_ MuI._1422_ vssd1 vssd1 vccd1 vccd1 MuI._1423_ sky130_fd_sc_hd__nor3_1
X_07724_ _00320_ _00325_ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__and2b_1
XMuI._6598_ MuI._0163_ MuI._0152_ MuI._0108_ vssd1 vssd1 vccd1 vccd1 MuI._2501_ sky130_fd_sc_hd__and3b_1
XFILLER_66_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5549_ MuI._1346_ MuI._1339_ vssd1 vssd1 vccd1 vccd1 MuI._1347_ sky130_fd_sc_hd__nor2_1
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07655_ _00268_ _00269_ _00270_ _00272_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__and4bb_1
XFILLER_198_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._429_ AuI.pe._393_ AuI.pe._394_ AuI.pe._395_ vssd1 vssd1 vccd1 vccd1 AuI.pe._396_
+ sky130_fd_sc_hd__and3_1
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10668__A _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _00188_ _00202_ _00203_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__nand3_1
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10387__B _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _01939_ _01941_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__nand3_1
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07042__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12801__A1 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09256_ _01866_ _01867_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__o21ai_2
XFILLER_194_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06881__A _04144_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ _00627_ _00625_ _00626_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__or3_1
XFILLER_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09187_ _02862_ _03993_ _01804_ _01802_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a31o_1
XANTENNA__07696__B _00307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _06622_ _05370_ _06489_ _00414_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__a22oi_2
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08069_ _00674_ _00675_ _00686_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__a21oi_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10100_ _02766_ _02769_ _02770_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__and4_1
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11080_ _03694_ _03828_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__xnor2_1
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10850__B _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _00955_ _00956_ _02700_ _01330_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07217__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11982_ _04796_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09432__A _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _03318_ _03490_ _02351_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__a21o_1
XFILLER_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1010_ AuI._0215_ AuI._0217_ AuI._0219_ AuI._0221_ AuI._0176_ AuI._0206_ vssd1
+ vssd1 vccd1 vccd1 AuI._0222_ sky130_fd_sc_hd__mux4_1
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10864_ _03460_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__and3_1
XANTENNA__13045__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _05421_ _05466_ _05468_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__or3_2
XFILLER_158_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ _03520_ _03521_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nor2_1
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07887__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _03024_ _05058_ _02744_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__a31o_1
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ _05309_ _05171_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__o21a_1
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._109_ FuI._052_ FuI._060_ FuI._064_ FuI.a_operand\[13\] vssd1 vssd1 vccd1 vccd1
+ FuI._003_ sky130_fd_sc_hd__o31a_1
XFILLER_172_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11416_ _00221_ _05456_ _04189_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a22o_1
X_12396_ _02324_ _02346_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__xor2_1
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4920_ MuI._0532_ MuI._0534_ vssd1 vssd1 vccd1 vccd1 MuI._0655_ sky130_fd_sc_hd__xor2_2
XANTENNA__12017__B _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11347_ _02980_ _00445_ _04907_ _02983_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a22o_1
XFILLER_180_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._780_ AuI.pe._003_ AuI.pe._040_ AuI.pe._118_ vssd1 vssd1 vccd1 vccd1 AuI.pe._321_
+ sky130_fd_sc_hd__or3_1
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4851_ MuI._0468_ MuI._0578_ vssd1 vssd1 vccd1 vccd1 MuI._0579_ sky130_fd_sc_hd__nor2_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output78_A net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11856__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _04038_ _04039_ _04040_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__a21o_1
XANTENNA__10760__B _03483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3802_ MuI._2900_ MuI._2901_ vssd1 vssd1 vccd1 vccd1 MuI._2902_ sky130_fd_sc_hd__nor2_1
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4782_ MuI.a_operand\[19\] MuI.a_operand\[18\] MuI.b_operand\[1\] MuI.b_operand\[0\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0503_ sky130_fd_sc_hd__and4_1
X_10229_ _05671_ _03507_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or2b_1
X_13017_ _05811_ _05812_ _05816_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__and3_1
XMuI._6521_ MuI._2406_ MuI._2405_ vssd1 vssd1 vccd1 vccd1 MuI._2416_ sky130_fd_sc_hd__and2b_1
XFILLER_94_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10334__A2 _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3733_ MuI._2824_ MuI._2832_ vssd1 vssd1 vccd1 vccd1 MuI._2833_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07127__A _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6111__A2 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6452_ MuI._2333_ MuI._2335_ vssd1 vssd1 vccd1 vccd1 MuI._2340_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3664_ MuI.a_operand\[14\] vssd1 vssd1 vccd1 vccd1 MuI._2660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5403_ MuI._2892_ MuI._2881_ MuI._0100_ MuI._3245_ vssd1 vssd1 vccd1 vccd1 MuI._1187_
+ sky130_fd_sc_hd__and4_1
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6383_ MuI._2257_ MuI._2262_ vssd1 vssd1 vccd1 vccd1 MuI._2265_ sky130_fd_sc_hd__or2_1
XMuI._3595_ MuI._1857_ MuI._1879_ vssd1 vssd1 vccd1 vccd1 MuI._1901_ sky130_fd_sc_hd__nand2_1
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5334_ MuI._1105_ MuI._1106_ MuI._1101_ MuI._1104_ vssd1 vssd1 vccd1 vccd1 MuI._1111_
+ sky130_fd_sc_hd__o211a_1
X_07440_ net119 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__buf_6
XAuI._1208_ AuI._0358_ AuI._0382_ AuI._0392_ AuI._0411_ vssd1 vssd1 vccd1 vccd1 AuI._0413_
+ sky130_fd_sc_hd__and4_1
XANTENNA__13036__A1 MuI.result\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0838__B_N net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5265_ MuI._2773_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._1035_ sky130_fd_sc_hd__nand2_1
XFILLER_195_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1139_ AuI._0256_ AuI._0343_ AuI._0345_ AuI._0346_ vssd1 vssd1 vccd1 vccd1 AuI._0348_
+ sky130_fd_sc_hd__a31o_1
X_07371_ _06670_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__and2b_1
XFILLER_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4216_ MuI._3091_ MuI._2898_ vssd1 vssd1 vccd1 vccd1 MuI._3316_ sky130_fd_sc_hd__nand2_1
X_09110_ _01724_ _01725_ _01726_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nand3_1
XANTENNA__11598__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5196_ MuI._2765_ MuI.a_operand\[9\] MuI._3402_ MuI._3396_ vssd1 vssd1 vccd1
+ vccd1 MuI._0959_ sky130_fd_sc_hd__and4_1
XANTENNA__07797__A _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4147_ MuI._3246_ vssd1 vssd1 vccd1 vccd1 MuI._3247_ sky130_fd_sc_hd__clkbuf_4
X_09041_ _01560_ _01562_ _01657_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__a211o_1
XANTENNA__10270__A1 _00691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4078_ MuI._3175_ MuI._3158_ vssd1 vssd1 vccd1 vccd1 MuI._3178_ sky130_fd_sc_hd__and2b_1
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1067__A1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._429__A AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09943_ _02603_ _02605_ _02592_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09715__A1 _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09715__B2 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09874_ _02118_ _02216_ _06437_ _04046_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__and4_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08140__B _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07682__D _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11522__A1 _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6719_ MuI._2389_ MuI._2633_ vssd1 vssd1 vccd1 vccd1 MuI._2634_ sky130_fd_sc_hd__and2_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07037__A _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5180__B MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08825_ _06495_ _06581_ _05101_ _02107_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22oi_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _06608_ _00272_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__nand2_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06876__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09252__A _01203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07707_ _00321_ _00324_ vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__xnor2_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6292__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _01303_ _01302_ _01301_ _01298_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__a211o_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07638_ _00254_ _00253_ _00148_ _00026_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__o211ai_2
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07569_ _00185_ _00184_ _00149_ _06659_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__o211a_1
XFILLER_167_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12786__B1 _05559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _01822_ _01814_ _01821_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._6169__A2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__A2 _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10580_ _03116_ _03113_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__and2b_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5058__D MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5636__A MuI._1438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10261__A1 AuI.result\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _01658_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__inv_2
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12250_ _04949_ _04950_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__a21oi_2
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12002__A2 _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _03956_ _03957_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__nand3_4
XANTENNA__11957__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _05007_ _03314_ _05009_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a31o_1
XFILLER_190_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11132_ _02983_ _02980_ _04789_ _00445_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nand4_2
XANTENNA__09427__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1490__B AuI._0542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6341__A2 MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10580__B _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ _03808_ _03799_ _03800_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and3_1
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1490_ AuI._0537_ AuI._0542_ vssd1 vssd1 vccd1 vccd1 AuI._0676_ sky130_fd_sc_hd__nor2_1
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08050__B _00519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10014_ _02665_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__xnor2_4
XFILLER_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09182__A2 _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4418__C MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06786__A _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3863__B1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4137__D MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _04780_ _04777_ _04779_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__nand3_1
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _03334_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__inv_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13018__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1368__D AuI._0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _03604_ _06605_ _06591_ _06434_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a22o_1
XFILLER_32_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ _03576_ _03577_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI._0850__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5050_ MuI._0796_ MuI._0797_ MuI._2966_ MuI._2319_ vssd1 vssd1 vccd1 vccd1 MuI._0798_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4001_ MuI._3098_ MuI._3099_ MuI._3090_ vssd1 vssd1 vccd1 vccd1 MuI._3101_ sky130_fd_sc_hd__a21o_1
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _02880_ _02885_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__nand2_1
XFILLER_201_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07410__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ _02711_ _05374_ _05375_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or3_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13497_ MuI.Exception _02739_ _02732_ AuI.Exception vssd1 vssd1 vccd1 vccd1 net101
+ sky130_fd_sc_hd__a22o_2
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5265__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12448_ _05291_ _05211_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__a21o_1
XFILLER_160_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5952_ MuI._1771_ MuI._1772_ MuI._1788_ MuI._1789_ vssd1 vssd1 vccd1 vccd1 MuI._1790_
+ sky130_fd_sc_hd__o211a_1
XANTENNA_MuI._4600__D MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11867__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _05146_ _05147_ _05226_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o211ai_4
XMuI._4903_ MuI._0447_ MuI._0446_ vssd1 vssd1 vccd1 vccd1 MuI._0637_ sky130_fd_sc_hd__and2b_1
XFILLER_126_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._832_ AuI.operand_a\[30\] AuI.pe._366_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[7\]
+ sky130_fd_sc_hd__xnor2_1
XMuI._5883_ MuI._1665_ MuI._1666_ vssd1 vssd1 vccd1 vccd1 MuI._1715_ sky130_fd_sc_hd__and2b_1
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._763_ AuI.pe.significand\[14\] AuI.pe._201_ AuI.pe._384_ AuI.pe._387_ AuI.pe._120_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._307_ sky130_fd_sc_hd__o2111a_1
XANTENNA_MuI._4343__A1 MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4834_ MuI._0556_ MuI._0558_ vssd1 vssd1 vccd1 vccd1 MuI._0561_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4343__B2 MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06940_ _04778_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__buf_6
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._694_ AuI.pe._386_ AuI.pe._238_ vssd1 vssd1 vccd1 vccd1 AuI.pe._241_ sky130_fd_sc_hd__xor2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4765_ MuI._0481_ MuI._0484_ vssd1 vssd1 vccd1 vccd1 MuI._0485_ sky130_fd_sc_hd__and2b_1
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06871_ _04035_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__buf_4
XMuI._6504_ MuI._2388_ MuI._2390_ MuI._2397_ vssd1 vssd1 vccd1 vccd1 MuI._2398_ sky130_fd_sc_hd__and3_1
XFILLER_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3716_ MuI._2812_ MuI._2815_ MuI._0867_ MuI._2363_ vssd1 vssd1 vccd1 vccd1 MuI._2816_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_83_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12400__A1_N _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ _01034_ _01226_ _01227_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__nand3_4
XFILLER_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4696_ MuI._0407_ MuI._0408_ vssd1 vssd1 vccd1 vccd1 MuI._0409_ sky130_fd_sc_hd__xnor2_1
X_09590_ _02223_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__xnor2_1
XMuI._6435_ MuI._2313_ MuI._2315_ MuI._2321_ vssd1 vssd1 vccd1 vccd1 MuI._2322_ sky130_fd_sc_hd__o21ba_1
XFILLER_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3647_ MuI.b_operand\[17\] vssd1 vssd1 vccd1 vccd1 MuI._2473_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09072__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ _00132_ _06433_ _04176_ _00133_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__a22oi_1
XANTENNA__08133__B1 _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6366_ MuI._1929_ MuI._1937_ vssd1 vssd1 vccd1 vccd1 MuI._2246_ sky130_fd_sc_hd__nand2_1
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3578_ MuI._1681_ MuI._1703_ vssd1 vssd1 vccd1 vccd1 MuI._1714_ sky130_fd_sc_hd__nand2_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _01082_ _01088_ _01089_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__a21bo_1
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5317_ MuI._0959_ MuI._0958_ MuI._0957_ vssd1 vssd1 vccd1 vccd1 MuI._1092_ sky130_fd_sc_hd__o21ai_1
XFILLER_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _00038_ _00039_ net121 _00040_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__and4b_1
XMuI._6297_ MuI._0746_ MuI._0790_ MuI._1153_ MuI._1032_ vssd1 vssd1 vccd1 vccd1 MuI._2170_
+ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3606__B1 MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5248_ MuI._0905_ MuI._0924_ MuI._0925_ vssd1 vssd1 vccd1 vccd1 MuI._1016_ sky130_fd_sc_hd__nand3_2
X_07354_ _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__B1 _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07320__A _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5179_ MuI._2583_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._0940_ sky130_fd_sc_hd__nand2_1
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07285_ _06583_ _04961_ _06584_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4360__A MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09024_ _01631_ _01632_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07947__B1 _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__C _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3704__A MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09926_ _02021_ _02027_ _02026_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a21o_1
XANTENNA__13496__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4885__A2 MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07990__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _02512_ _02504_ _02511_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__or3b_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08372__B1 _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08808_ _01424_ _01425_ _00444_ _03873_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and4bb_1
XFILLER_65_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _02436_ _02437_ _02429_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nor3b_2
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _01354_ _01356_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__nor2_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _04512_ _04549_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__or3_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09710__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10701_ _06598_ _06599_ _06476_ _06489_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__and4_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _04291_ _04293_ _04475_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a211o_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13420_ _02823_ _02824_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nor2_1
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ _03143_ _03146_ _03144_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12223__A2 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5366__A MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13351_ _03561_ _05724_ _02742_ _02943_ _05671_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a32o_1
X_10563_ _03097_ _03095_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._6011__A1 MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0990_ AuI._0175_ AuI._0199_ AuI._0200_ AuI._0201_ vssd1 vssd1 vccd1 vccd1 AuI._0202_
+ sky130_fd_sc_hd__and4_1
XFILLER_195_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6011__B2 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10785__A2 _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _04975_ _05076_ _05114_ _05115_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a211oi_2
XFILLER_182_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ _01147_ _01146_ _04714_ _04789_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and4_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _06047_ _06049_ _06130_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__and3_1
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _05068_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__nand2_1
XFILLER_170_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11734__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__B1 _00555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1611_ AuI._0779_ AuI._0780_ vssd1 vssd1 vccd1 vccd1 AuI._0781_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11734__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _04993_ _04995_ _04864_ _04868_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__o211a_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11115_ _00678_ _00047_ _00048_ _06434_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a22o_1
XAuI._1542_ AuI._0723_ AuI._0659_ vssd1 vssd1 vccd1 vccd1 AuI._0724_ sky130_fd_sc_hd__xor2_1
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12095_ _03324_ _05391_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XANTENNA__13487__A1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11046_ _03789_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__nand3_1
XANTENNA__08211__D net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1473_ AuI._0382_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0659_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6078__A1 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5251__D MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4550_ MuI._0243_ MuI._0247_ vssd1 vssd1 vccd1 vccd1 MuI._0248_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__A2 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__A _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13239__A1 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3501_ MuI.b_operand\[20\] vssd1 vssd1 vccd1 vccd1 MuI._0867_ sky130_fd_sc_hd__buf_2
XANTENNA__13239__B2 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4481_ MuI._0169_ MuI._0170_ MuI._0171_ vssd1 vssd1 vccd1 vccd1 MuI._0172_ sky130_fd_sc_hd__o21ba_1
XFILLER_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6220_ MuI._0867_ MuI._2849_ MuI._2051_ MuI._2052_ vssd1 vssd1 vccd1 vccd1 MuI._2085_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ _05804_ _05807_ _05805_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__o21ba_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3432_ MuI.a_operand\[29\] MuI.b_operand\[29\] vssd1 vssd1 vccd1 vccd1 MuI._0108_
+ sky130_fd_sc_hd__nand2_1
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07124__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07469__A2 _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _04761_ _04762_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__a21oi_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6151_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._2649_ vssd1 vssd1 vccd1
+ vccd1 MuI._2009_ sky130_fd_sc_hd__o31a_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._5102_ MuI.a_operand\[11\] MuI.a_operand\[10\] MuI._0017_ MuI._0018_ vssd1 vssd1
+ vccd1 vccd1 MuI._0855_ sky130_fd_sc_hd__and4_1
X_11879_ _04687_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__and3_1
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6082_ MuI._1472_ MuI._1802_ MuI._2843_ MuI._1307_ vssd1 vssd1 vccd1 vccd1 MuI._1933_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_177_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08881__D net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5033_ MuI._0776_ MuI._0777_ vssd1 vssd1 vccd1 vccd1 MuI._0780_ sky130_fd_sc_hd__nor2_1
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4180__A MuI._3278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4831__A1_N MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5707__C MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__A _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ _04262_ _06067_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__and2_1
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3508__B MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07929__B1 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5935_ MuI._1735_ MuI._1753_ vssd1 vssd1 vccd1 vccd1 MuI._1772_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._6305__A2 MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._815_ AuI.pe._367_ AuI.pe._368_ AuI.pe._369_ AuI.pe._372_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._354_ sky130_fd_sc_hd__or4_1
XANTENNA__12205__B _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5866_ MuI._1687_ MuI._1688_ MuI._1695_ vssd1 vssd1 vccd1 vccd1 MuI._1696_ sky130_fd_sc_hd__and3_1
XFILLER_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07972_ _00304_ _00589_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__nor2_1
XMuI._4817_ MuI._0539_ MuI._0540_ MuI._0541_ vssd1 vssd1 vccd1 vccd1 MuI._0542_ sky130_fd_sc_hd__a21boi_1
XAuI.pe._746_ AuI.pe.significand\[21\] AuI.pe._270_ vssd1 vssd1 vccd1 vccd1 AuI.pe._291_
+ sky130_fd_sc_hd__or2_1
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09711_ _02353_ _02354_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__xor2_1
XMuI._5797_ MuI._1612_ MuI._1613_ MuI._1619_ vssd1 vssd1 vccd1 vccd1 MuI._1620_ sky130_fd_sc_hd__nand3_1
X_06923_ _04596_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._677_ AuI.pe._062_ AuI.pe._197_ AuI.pe._010_ vssd1 vssd1 vccd1 vccd1 AuI.pe._225_
+ sky130_fd_sc_hd__and3_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4748_ MuI.a_operand\[14\] MuI.a_operand\[13\] MuI._2866_ MuI._2868_ vssd1 vssd1
+ vccd1 vccd1 MuI._0466_ sky130_fd_sc_hd__and4_1
XFILLER_28_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _02278_ _02279_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o21ba_1
XFILLER_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13317__A _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ _03852_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[31\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__12221__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__A2 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4679_ MuI._0160_ MuI._0161_ vssd1 vssd1 vccd1 vccd1 MuI._0390_ sky130_fd_sc_hd__nor2_1
X_06785_ _02042_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__clkbuf_2
X_09573_ _02189_ _02190_ _02203_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a21o_1
XFILLER_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6418_ MuI._2289_ MuI._2302_ vssd1 vssd1 vccd1 vccd1 MuI._2303_ sky130_fd_sc_hd__nand2_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08524_ _01138_ _01139_ _01141_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__o21ai_1
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4074__B MuI._3171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__B _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6349_ MuI._2213_ MuI._2226_ vssd1 vssd1 vccd1 vccd1 MuI._2227_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ _00029_ _00072_ _00083_ _00028_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__a22oi_2
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07406_ _06676_ _06677_ _00023_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__o21a_1
X_08386_ _00832_ _00824_ _00831_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__nand3_1
XFILLER_196_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._090_ FuI._050_ vssd1 vssd1 vccd1 vccd1 FuI._052_ sky130_fd_sc_hd__buf_2
XANTENNA__07050__A _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ _06617_ _06618_ _06636_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__nand3_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4521__C MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A2 _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _06560_ _06568_ _06563_ _06566_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__a22o_1
XFILLER_164_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _01618_ _01621_ _01590_ _01591_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a211o_1
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07199_ net109 vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__buf_4
XFILLER_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11716__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11716__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07396__A1 _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__D _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5504__B1 MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13469__A1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09909_ _02518_ _02525_ _02545_ _02524_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__o22ai_1
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3530__A2 MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12920_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__D _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07225__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12851_ _05694_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__xnor2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11802_ _04440_ _04442_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__nor2_1
XFILLER_199_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _05555_ _05557_ _05658_ _05659_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a211oi_4
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _04530_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nand2_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4243__B1 MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11664_ _04457_ _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nand3_1
XANTENNA__07871__A2 _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ _02817_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nand2_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11404__B1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ _03290_ _03292_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nor2_1
XFILLER_195_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11595_ _04219_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__inv_2
XFILLER_167_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11955__A1 _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11955__B2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334_ _06185_ _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nand2_1
X_10546_ _03252_ _03253_ _03244_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a21o_1
XAuI._0973_ AuI._0164_ AuI._0169_ AuI._0184_ vssd1 vssd1 vccd1 vccd1 AuI._0185_ sky130_fd_sc_hd__and3_1
XFILLER_183_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ _06017_ _06108_ _06111_ _06109_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__o22a_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10477_ _03139_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__xor2_2
XFILLER_170_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3981_ MuI._3071_ MuI._3080_ vssd1 vssd1 vccd1 vccd1 MuI._3081_ sky130_fd_sc_hd__nand2_1
X_12216_ _03335_ _05456_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nand2_2
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13196_ _03507_ _05992_ _06039_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__a21oi_1
XMuI._5720_ MuI._1532_ MuI._1533_ MuI._1524_ vssd1 vssd1 vccd1 vccd1 MuI._1535_ sky130_fd_sc_hd__a21o_1
XFILLER_124_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _04975_ _04976_ _04956_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5262__C MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._600_ AuI.pe._125_ AuI.pe._041_ AuI.pe._119_ AuI.pe.significand\[2\] AuI.pe._153_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._154_ sky130_fd_sc_hd__a221o_1
XMuI._5651_ MuI._1062_ MuI._1172_ MuI._1178_ vssd1 vssd1 vccd1 vccd1 MuI._1459_ sky130_fd_sc_hd__nor3_1
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1525_ AuI._0599_ AuI._0692_ vssd1 vssd1 vccd1 vccd1 AuI._0709_ sky130_fd_sc_hd__and2_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._531_ AuI.pe._089_ AuI.pe._026_ AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 AuI.pe._090_
+ sky130_fd_sc_hd__a21o_1
XFILLER_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12078_ _04828_ _04829_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or2_1
XMuI._4602_ MuI._0304_ vssd1 vssd1 vccd1 vccd1 MuI._0305_ sky130_fd_sc_hd__buf_4
XFILLER_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5582_ MuI._1353_ MuI._1350_ MuI._1352_ vssd1 vssd1 vccd1 vccd1 MuI._1383_ sky130_fd_sc_hd__or3_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11029_ _03617_ _03619_ _03772_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a211oi_4
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1456_ AuI._0462_ AuI._0467_ AuI._0641_ vssd1 vssd1 vccd1 vccd1 AuI._0642_ sky130_fd_sc_hd__o21a_1
XAuI.pe._462_ AuI.pe._024_ AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 AuI.pe._027_ sky130_fd_sc_hd__and2_1
XFILLER_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4533_ MuI.b_operand\[19\] MuI._2811_ MuI._2829_ MuI._0228_ vssd1 vssd1 vccd1
+ vccd1 MuI._0230_ sky130_fd_sc_hd__and4_1
XFILLER_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07135__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3809__B1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1387_ AuI._0257_ AuI._0575_ AuI._0576_ AuI._0577_ vssd1 vssd1 vccd1 vccd1 AuI._0578_
+ sky130_fd_sc_hd__nand4_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4464_ MuI._0023_ MuI._0153_ vssd1 vssd1 vccd1 vccd1 MuI._0154_ sky130_fd_sc_hd__nor2_1
XANTENNA_AuI.pe._667__A2 AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6203_ MuI._1887_ MuI._2065_ MuI._2851_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._2067_
+ sky130_fd_sc_hd__o211a_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06974__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4395_ MuI._2796_ MuI._2786_ vssd1 vssd1 vccd1 vccd1 MuI._0078_ sky130_fd_sc_hd__nand2_1
XANTENNA__09300__A2 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6223__A1 MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10496__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6134_ MuI._1985_ MuI._1988_ vssd1 vssd1 vccd1 vccd1 MuI._1991_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._6223__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08240_ _00851_ _00856_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__xor2_1
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6065_ MuI._1911_ MuI._1914_ vssd1 vssd1 vccd1 vccd1 MuI._1915_ sky130_fd_sc_hd__or2b_1
XANTENNA__13396__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08171_ net29 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_4
XFILLER_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09064__A1 _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09064__B2 _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5016_ MuI._0585_ MuI._0759_ MuI._0758_ MuI._0754_ vssd1 vssd1 vccd1 vccd1 MuI._0761_
+ sky130_fd_sc_hd__a211oi_1
XANTENNA_MuI._4341__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07122_ _05917_ _06056_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__and2_1
XFILLER_174_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07614__A2 _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5156__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07053_ _05992_ _02042_ _02151_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__and3_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 ALU_Output[9] sky130_fd_sc_hd__buf_2
XFILLER_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12216__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5918_ MuI._1737_ MuI._1752_ vssd1 vssd1 vccd1 vccd1 MuI._1753_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5849_ MuI._0712_ MuI._1676_ vssd1 vssd1 vccd1 vccd1 MuI._1677_ sky130_fd_sc_hd__nor2_1
X_07955_ _00062_ _00085_ _04585_ _00063_ vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a22oi_2
XANTENNA_MuI._4170__C1 MuI._0515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._729_ AuI.pe._273_ AuI.pe._375_ AuI.pe._376_ vssd1 vssd1 vccd1 vccd1 AuI.pe._274_
+ sky130_fd_sc_hd__nor3_1
XFILLER_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06906_ _04413_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[7\] sky130_fd_sc_hd__clkbuf_2
XANTENNA__11493__C _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ _06441_ _06448_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__and2_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07045__A _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _02258_ _02261_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__nand3_1
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06837_ _03669_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__buf_2
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _02139_ _02141_ _02142_ _02087_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__o22ai_1
XFILLER_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06768_ _02927_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[15\] sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06884__A _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08507_ _01108_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _06548_ _04434_ _00098_ _02291_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22oi_1
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06699_ net116 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__clkbuf_4
XFILLER_169_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08438_ _01038_ _01043_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__nand2_1
XFILLER_211_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._142_ FuI._004_ net148 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[13\] sky130_fd_sc_hd__dlxtn_1
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13387__B1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11014__B _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08369_ _00970_ _00985_ _00984_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__a21o_1
XFILLER_165_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFuI._073_ FuI.a_operand\[23\] FuI._035_ FuI._040_ FuI.a_operand\[1\] vssd1 vssd1
+ vccd1 vccd1 FuI._010_ sky130_fd_sc_hd__o211a_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _00781_ _00797_ _03096_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__o21a_1
XFILLER_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08604__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _03021_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nor2_1
XANTENNA__12126__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10262_ _02216_ _04004_ _02724_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__o21a_1
X_13050_ _05944_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nor2_1
XFILLER_180_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _04819_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__xor2_1
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10193_ _00789_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__inv_2
XFILLER_132_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09435__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1310_ AuI._0437_ AuI._0502_ AuI._0505_ AuI._0506_ vssd1 vssd1 vccd1 vccd1 AuI._0508_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0917__A0 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _05787_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor2_1
XAuI._1241_ net36 net68 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0444_ sky130_fd_sc_hd__mux2_1
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11873__B1 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12796__A _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1172_ AuI._0256_ AuI._0377_ AuI._0378_ vssd1 vssd1 vccd1 vccd1 AuI._0379_ sky130_fd_sc_hd__nand3_1
X_12834_ _06442_ _03051_ _03071_ _06444_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__a22oi_1
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06794__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10428__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__A2 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12765_ _05519_ _05521_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a21o_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6205__A1 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A2 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4180_ MuI._3278_ MuI._3279_ vssd1 vssd1 vccd1 vccd1 MuI._3280_ sky130_fd_sc_hd__xor2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11716_ _00046_ _00382_ _00163_ _00049_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a22o_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12696_ _05346_ _05480_ _05481_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__o21a_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11647_ _04438_ _04439_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__xnor2_4
XFILLER_156_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 a_operand[17] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_6
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput24 a_operand[27] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_4
Xinput35 a_operand[8] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 b_operand[18] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_6
X_11578_ _04050_ _04246_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__nor2_1
XFILLER_183_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 b_operand[28] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_4
XFILLER_171_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput68 b_operand[9] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_4
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10600__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13317_ _03680_ _05981_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nand2_1
X_10529_ _03226_ _03234_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__nand3_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0956_ AuI._0165_ AuI._0167_ AuI._0117_ vssd1 vssd1 vccd1 vccd1 AuI._0168_ sky130_fd_sc_hd__a21o_1
XFILLER_155_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6821_ MuI._2741_ vssd1 vssd1 vccd1 vccd1 MuI.result\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13248_ _06100_ _06143_ _06149_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__or4b_4
XAuI._0887_ net56 vssd1 vssd1 vccd1 vccd1 AuI._0107_ sky130_fd_sc_hd__inv_2
XFILLER_130_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11156__A2 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3964_ MuI._3062_ MuI._3063_ vssd1 vssd1 vccd1 vccd1 MuI._3064_ sky130_fd_sc_hd__xor2_1
XMuI._6752_ MuI._2482_ MuI._2505_ MuI._2668_ MuI._2669_ vssd1 vssd1 vccd1 vccd1 MuI._2670_
+ sky130_fd_sc_hd__o31ai_1
XFILLER_124_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11875__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _02708_ _02841_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__nor2_1
XFILLER_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06969__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5703_ MuI._1512_ MuI._1513_ MuI._1514_ vssd1 vssd1 vccd1 vccd1 MuI._1517_ sky130_fd_sc_hd__o21ai_1
XMuI._6683_ MuI._2590_ MuI._2593_ MuI._2485_ vssd1 vssd1 vccd1 vccd1 MuI._2595_ sky130_fd_sc_hd__mux2_1
XFILLER_112_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3895_ MuI._2972_ MuI._2988_ MuI._2989_ MuI._2994_ vssd1 vssd1 vccd1 vccd1 MuI._2995_
+ sky130_fd_sc_hd__a31o_1
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4298__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5634_ MuI._1418_ MuI._1440_ vssd1 vssd1 vccd1 vccd1 MuI._1441_ sky130_fd_sc_hd__nor2_1
XANTENNA__13302__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1508_ AuI._0608_ AuI._0612_ AuI._0693_ vssd1 vssd1 vccd1 vccd1 AuI._0694_ sky130_fd_sc_hd__mux2_1
X_07740_ _00356_ _00357_ vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__nor2_1
XFILLER_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._514_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._074_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4617__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5565_ MuI._1360_ MuI._1364_ vssd1 vssd1 vccd1 vccd1 MuI._1365_ sky130_fd_sc_hd__and2b_1
XFILLER_65_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10667__A1 _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1439_ AuI._0515_ AuI._0519_ vssd1 vssd1 vccd1 vccd1 AuI._0625_ sky130_fd_sc_hd__xor2_1
X_07671_ _03432_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__buf_4
XMuI._4516_ MuI._2649_ MuI._2773_ MuI._2786_ MuI._2704_ vssd1 vssd1 vccd1 vccd1 MuI._0211_
+ sky130_fd_sc_hd__a22oi_2
XAuI.pe._445_ AuI.pe.significand\[4\] AuI.pe._388_ AuI.pe._009_ AuI.pe._011_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._012_ sky130_fd_sc_hd__and4_1
XFILLER_93_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09410_ _01952_ _01954_ _01953_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a21oi_1
XMuI._5496_ MuI._1242_ MuI._1287_ MuI._1183_ MuI._1235_ vssd1 vssd1 vccd1 vccd1 MuI._1289_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_198_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4447_ MuI._3368_ MuI._3373_ MuI._3369_ vssd1 vssd1 vccd1 vccd1 MuI._0135_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09080__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _01882_ _01883_ _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__and3_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4378_ MuI._0058_ MuI._0056_ vssd1 vssd1 vccd1 vccd1 MuI._0060_ sky130_fd_sc_hd__xnor2_1
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11092__B2 _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _06564_ _00082_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand2_1
XFILLER_194_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6117_ MuI._0559_ MuI._0768_ MuI._2693_ MuI._2638_ vssd1 vssd1 vccd1 vccd1 MuI._1972_
+ sky130_fd_sc_hd__and4_1
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08223_ _02485_ _06584_ _05112_ _06565_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a22oi_2
XFILLER_194_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6048_ MuI._1032_ MuI._2800_ MuI._2919_ MuI._0790_ vssd1 vssd1 vccd1 vccd1 MuI._1896_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _00383_ _00386_ _00384_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__o21bai_1
XANTENNA__11395__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _06416_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[21\] sky130_fd_sc_hd__clkbuf_1
XFILLER_174_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08085_ _00692_ _00701_ _00702_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__and3_1
XFILLER_162_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07036_ net128 vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06879__A _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0927__B AuI._0138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07220__B1 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08987_ _01602_ _01603_ _01604_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nand3_2
XFILLER_130_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3497__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _02765_ _04854_ _00555_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11855__B1 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _00279_ _00074_ _00090_ _00278_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _02199_ _02198_ _02197_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _03609_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a21o_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08981__A2_N _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _02168_ _02169_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__and2_1
XANTENNA_AuI.pe._500__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09276__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1324__B1 AuI._0519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ _05408_ _05409_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__and3_1
XFILLER_169_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11501_ _04271_ _04281_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__and3_1
XFILLER_200_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4749__B2 MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ _05222_ _05224_ _05335_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o211a_1
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._125_ net104 FuI._026_ FuI.a_operand\[20\] net105 vssd1 vssd1 vccd1 vccd1 FuI._011_
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1493__B AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ _00132_ _05316_ _05380_ _00133_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__a22oi_1
XFILLER_165_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__A1 _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__B2 _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0810_ AuI._0025_ net114 vssd1 vssd1 vccd1 vccd1 AuI._0030_ sky130_fd_sc_hd__and2_1
X_11363_ _04131_ _04132_ _04113_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__a21o_1
XFILLER_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5174__A1 MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ _05467_ _02941_ _02782_ _03306_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__o22ai_1
XANTENNA_MuI._5174__B2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10314_ _00725_ _00745_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__nor2_1
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11294_ _00444_ _05391_ _04056_ _04058_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__nand4_1
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13033_ _02779_ _05927_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_152_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10245_ _06045_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09200__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09200__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06789__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _02854_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__nand2_2
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3680_ MuI._2759_ MuI._2778_ MuI._2779_ vssd1 vssd1 vccd1 vccd1 MuI._2780_ sky130_fd_sc_hd__or3_1
XFILLER_93_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12099__B1 _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5540__C MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5350_ MuI._1126_ MuI._1127_ vssd1 vssd1 vccd1 vccd1 MuI._1128_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1224_ net35 net67 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0428_ sky130_fd_sc_hd__mux2_1
XFILLER_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4301_ MuI._0570_ MuI._3269_ MuI._3399_ MuI._3400_ vssd1 vssd1 vccd1 vccd1 MuI._3401_
+ sky130_fd_sc_hd__a31o_1
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5281_ MuI._0924_ MuI._1016_ MuI._1050_ MuI._1051_ vssd1 vssd1 vccd1 vccd1 MuI._1052_
+ sky130_fd_sc_hd__a211oi_4
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07413__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1155_ AuI._0256_ AuI._0359_ AuI._0360_ AuI._0361_ vssd1 vssd1 vccd1 vccd1 AuI._0363_
+ sky130_fd_sc_hd__a31o_1
X_12817_ _05604_ _05607_ _05603_ _05602_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09267__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09267__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4232_ MuI._3329_ MuI._3331_ vssd1 vssd1 vccd1 vccd1 MuI._3332_ sky130_fd_sc_hd__and2b_1
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _05620_ _05621_ _05614_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a21o_1
XAuI._1086_ AuI._0261_ AuI._0289_ AuI._0296_ vssd1 vssd1 vccd1 vccd1 AuI._0297_ sky130_fd_sc_hd__and3_1
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12810__A2 _05959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4163_ MuI.a_operand\[22\] MuI._3262_ vssd1 vssd1 vccd1 vccd1 MuI._3263_ sky130_fd_sc_hd__and2_1
XFILLER_188_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ _05547_ _05548_ _05419_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4094_ MuI._2077_ MuI._2898_ MuI._3193_ MuI._3191_ vssd1 vssd1 vccd1 vccd1 MuI._3194_
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__B _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08242__A2 _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._558__B2 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0939_ AuI._0097_ AuI._0147_ AuI._0149_ vssd1 vssd1 vccd1 vccd1 AuI._0151_ sky130_fd_sc_hd__nand3_1
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6804_ MuI._2653_ MuI._2676_ MuI._2656_ vssd1 vssd1 vccd1 vccd1 MuI._2728_ sky130_fd_sc_hd__a21o_1
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3715__A2 MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _01512_ _01513_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a21o_1
XFILLER_98_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4996_ MuI._0636_ MuI._0421_ MuI._0644_ MuI._0738_ vssd1 vssd1 vccd1 vccd1 MuI._0739_
+ sky130_fd_sc_hd__a31oi_4
X_09890_ _02450_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06699__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6735_ MuI._2424_ MuI._2651_ vssd1 vssd1 vccd1 vccd1 MuI._2652_ sky130_fd_sc_hd__xnor2_1
XMuI._3947_ MuI._3043_ MuI._3044_ MuI._3045_ vssd1 vssd1 vccd1 vccd1 MuI._3047_ sky130_fd_sc_hd__a21o_1
X_08841_ _06534_ _06491_ _06580_ _06581_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__nand4_1
XFILLER_98_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3532__A MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3878_ MuI._2973_ MuI._2974_ MuI._2977_ vssd1 vssd1 vccd1 vccd1 MuI._2978_ sky130_fd_sc_hd__or3_1
XMuI._6666_ MuI._2568_ MuI._2571_ MuI._2575_ vssd1 vssd1 vccd1 vccd1 MuI._2576_ sky130_fd_sc_hd__and3_1
XFILLER_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _00028_ _00029_ _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__and4_1
XFILLER_100_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12629__A2 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5617_ MuI._1420_ MuI._1415_ MuI._1418_ vssd1 vssd1 vccd1 vccd1 MuI._1422_ sky130_fd_sc_hd__nor3_1
XANTENNA__09803__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _00328_ vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XMuI._6597_ MuI._0207_ MuI._2498_ MuI._2499_ vssd1 vssd1 vccd1 vccd1 MuI._2500_ sky130_fd_sc_hd__a21o_1
XANTENNA__11837__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5548_ MuI._1336_ MuI._1337_ MuI._1338_ vssd1 vssd1 vccd1 vccd1 MuI._1346_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07654_ _00271_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__buf_4
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._428_ AuI.pe._367_ AuI.pe._368_ AuI.pe._369_ AuI.pe._372_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._395_ sky130_fd_sc_hd__nor4_4
XANTENNA__10668__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5459__A MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5479_ MuI._1202_ MuI._1212_ MuI._1213_ vssd1 vssd1 vccd1 vccd1 MuI._1270_ sky130_fd_sc_hd__and3_1
XFILLER_198_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07323__A _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__C _01266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07585_ _00195_ _00196_ _00201_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__a21o_1
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _01926_ _01938_ _01937_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a21o_1
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12801__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._450__A AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _01868_ _01872_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10684__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _00822_ _00823_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12014__B1 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ _01802_ _01803_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._5194__A MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08137_ _00753_ _00754_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ _00684_ _00685_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__xor2_1
XANTENNA_AuI._0832__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07019_ _05627_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__clkbuf_4
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _01200_ _01320_ _01326_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4667__B1 MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11981_ _04796_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__and3_1
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _02564_ _03314_ _03668_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__and3b_1
XANTENNA__09432__B _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1488__B AuI._0542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07233__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4273__A MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _03591_ _03592_ _03393_ _03413_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__o211a_1
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13045__A2 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6191__C MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11056__A1 _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ _05464_ _05465_ _05422_ _05326_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a211oi_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3642__A1 MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _00506_ _03604_ _04445_ _00085_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__and4_1
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12533_ _05058_ _02727_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__nor2_1
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07887__B _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12464_ _05310_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__xor2_1
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._108_ FuI._037_ FuI._056_ FuI._058_ vssd1 vssd1 vccd1 vccd1 FuI._064_ sky130_fd_sc_hd__and3b_1
XFILLER_138_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _02905_ _02959_ _03051_ _03071_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nand4_1
X_12395_ _05240_ _05243_ _03133_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__o21a_1
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__A_N _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07432__B1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11346_ _03962_ _03965_ _03963_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__o21bai_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0848__A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4850_ MuI._2451_ MuI._0168_ MuI._0466_ MuI._0467_ vssd1 vssd1 vccd1 vccd1 MuI._0578_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11856__C _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _04038_ _04039_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nand3_1
XFILLER_140_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3801_ MuI._0779_ MuI._2874_ MuI._2876_ MuI._2894_ vssd1 vssd1 vccd1 vccd1 MuI._2901_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__09185__B1 _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4781_ MuI._0422_ MuI._0500_ MuI._0501_ vssd1 vssd1 vccd1 vccd1 MuI._0502_ sky130_fd_sc_hd__a21o_1
X_13016_ _05826_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__xnor2_1
X_10228_ _02836_ _02838_ _02834_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__o21a_1
XFILLER_79_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3732_ MuI._2828_ MuI._2831_ vssd1 vssd1 vccd1 vccd1 MuI._2832_ sky130_fd_sc_hd__xnor2_1
XMuI._6520_ MuI._2264_ MuI._2399_ MuI._2414_ vssd1 vssd1 vccd1 vccd1 MuI._2415_ sky130_fd_sc_hd__or3b_1
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__nor2_2
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3663_ MuI._2638_ vssd1 vssd1 vccd1 vccd1 MuI._2649_ sky130_fd_sc_hd__buf_2
XFILLER_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6451_ MuI._2337_ MuI._2338_ vssd1 vssd1 vccd1 vccd1 MuI._2339_ sky130_fd_sc_hd__or2_1
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11819__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12062__A1_N _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5402_ MuI._1137_ MuI._1136_ MuI._1128_ vssd1 vssd1 vccd1 vccd1 MuI._1185_ sky130_fd_sc_hd__a21o_1
XMuI._6382_ MuI._2257_ MuI._2262_ vssd1 vssd1 vccd1 vccd1 MuI._2263_ sky130_fd_sc_hd__nand2_1
XFILLER_63_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3594_ MuI._1329_ MuI._1285_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._1890_ sky130_fd_sc_hd__and3b_1
XFILLER_208_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5333_ MuI._1067_ MuI._1083_ vssd1 vssd1 vccd1 vccd1 MuI._1110_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07143__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1207_ AuI._0367_ AuI._0382_ AuI._0392_ AuI._0411_ vssd1 vssd1 vccd1 vccd1 AuI._0412_
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._4183__A MuI._3160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5264_ MuI._1031_ MuI._1033_ vssd1 vssd1 vccd1 vccd1 MuI._1034_ sky130_fd_sc_hd__nor2_1
XFuI._130__136 vssd1 vssd1 vccd1 vccd1 FuI._130__136/HI net136 sky130_fd_sc_hd__conb_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1138_ AuI._0256_ AuI._0343_ AuI._0345_ AuI._0346_ vssd1 vssd1 vccd1 vccd1 AuI._0347_
+ sky130_fd_sc_hd__and4_1
XFILLER_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ _06668_ _06669_ _06662_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a21o_1
XANTENNA__06982__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4215_ MuI._3308_ MuI._3312_ MuI._3314_ vssd1 vssd1 vccd1 vccd1 MuI._3315_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__A2 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5195_ MuI._2785_ MuI._3262_ MuI._0020_ MuI._2790_ vssd1 vssd1 vccd1 vccd1 MuI._0958_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07797__B _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1069_ AuI._0223_ AuI._0199_ AuI._0200_ AuI._0279_ vssd1 vssd1 vccd1 vccd1 AuI._0280_
+ sky130_fd_sc_hd__and4_1
XMuI._4146_ MuI._3245_ vssd1 vssd1 vccd1 vccd1 MuI._3246_ sky130_fd_sc_hd__clkbuf_4
X_09040_ _01650_ _01651_ _01656_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__and3_1
XFILLER_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3527__A MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4077_ MuI._2418_ MuI._2958_ vssd1 vssd1 vccd1 vccd1 MuI._3177_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5742__A MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _02034_ _02591_ _02590_ _02588_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__o211a_1
XANTENNA__09715__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4979_ MuI._0624_ MuI._0715_ vssd1 vssd1 vccd1 vccd1 MuI._0720_ sky130_fd_sc_hd__nor2_1
X_09873_ _02503_ _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4358__A MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07726__A1 _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6718_ MuI._2306_ MuI._2628_ vssd1 vssd1 vccd1 vccd1 MuI._2633_ sky130_fd_sc_hd__or2b_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07726__B2 _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11522__A2 _04303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _06460_ net133 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__nand2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__B1 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._445__A AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6649_ MuI._2553_ MuI._2555_ MuI._2556_ vssd1 vssd1 vccd1 vccd1 MuI._2557_ sky130_fd_sc_hd__or3_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08755_ _01371_ _01369_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__xnor2_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _00322_ _00323_ vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__and2b_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09252__B _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08686_ _01298_ _01301_ _01302_ _01303_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__o211ai_4
XFILLER_199_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6292__B MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07053__A _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1_N _03913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _00026_ _00148_ _00253_ _00254_ vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__a211o_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06892__A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _06659_ _00149_ _00184_ _00185_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__a211oi_4
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09307_ _01809_ _01838_ _01839_ _01837_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__o22a_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07499_ _00112_ _00114_ _00113_ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__a21o_1
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10261__A2 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _01854_ _01853_ _01852_ _01631_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a211oi_1
XFILLER_194_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09169_ _02582_ _02647_ _00266_ _00592_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._5355__C MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _03750_ _03749_ _03748_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12180_ _02808_ _02724_ _05010_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a211o_1
XANTENNA__11957__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _03443_ _06612_ _04843_ _00290_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__a22o_1
XANTENNA__09427__B _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12134__A _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _03799_ _03800_ _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _01319_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__nor2_2
XFILLER_0_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10721__B1 _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A a_operand[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4418__D MuI._0101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3900__A MuI.b_operand\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3863__A1 MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _04777_ _04779_ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._3863__B2 MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10036__B_N net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10915_ _03513_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__xnor2_4
XFILLER_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13018__A2 _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895_ _06434_ _03604_ _06605_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__and3_1
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10846_ _00270_ _04789_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__nand2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4000_ MuI._3090_ MuI._3098_ MuI._3099_ vssd1 vssd1 vccd1 vccd1 MuI._3100_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4731__A MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ _02563_ _03315_ _03316_ _03502_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__a31o_4
XFILLER_197_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11213__A _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _05363_ _05373_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and2_1
XFILLER_158_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13496_ _04161_ _02813_ _06409_ _02739_ MuI.Overflow vssd1 vssd1 vccd1 vccd1 net102
+ sky130_fd_sc_hd__a32o_4
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12529__A1 _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__xor2_1
XFILLER_173_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output90_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5951_ MuI._1787_ MuI._1786_ MuI._1782_ vssd1 vssd1 vccd1 vccd1 MuI._1789_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._4591__A2 MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11867__B _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ _05224_ _05225_ _05180_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__o21ai_2
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._831_ AuI.pe._360_ AuI.pe._362_ AuI.pe._364_ AuI.operand_a\[29\] vssd1 vssd1
+ vccd1 vccd1 AuI.pe._366_ sky130_fd_sc_hd__a211o_1
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4902_ MuI._0625_ MuI._0420_ vssd1 vssd1 vccd1 vccd1 MuI._0635_ sky130_fd_sc_hd__nand2_1
XFILLER_153_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5882_ MuI._1647_ MuI._1710_ vssd1 vssd1 vccd1 vccd1 MuI._1713_ sky130_fd_sc_hd__nand2_1
XFILLER_141_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _03879_ _03898_ _03899_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__and3_1
XANTENNA__12044__A _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08241__B _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._762_ AuI.pe.significand\[21\] AuI.pe._025_ AuI.pe.significand\[22\] AuI.pe.significand\[24\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._306_ sky130_fd_sc_hd__o211a_1
XANTENNA__10960__B1 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4343__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4833_ MuI._0556_ MuI._0558_ vssd1 vssd1 vccd1 vccd1 MuI._0560_ sky130_fd_sc_hd__and2b_1
XFILLER_141_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07138__A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._693_ AuI.pe._227_ AuI.pe._237_ AuI.pe._240_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[18\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__08905__B1 _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4764_ MuI._0331_ MuI._0483_ vssd1 vssd1 vccd1 vccd1 MuI._0484_ sky130_fd_sc_hd__nor2_1
X_06870_ net127 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06977__A _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6503_ MuI._2392_ MuI._2395_ MuI._2367_ vssd1 vssd1 vccd1 vccd1 MuI._2397_ sky130_fd_sc_hd__a21o_1
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3715_ MuI._2813_ MuI._2773_ MuI._2786_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._2815_
+ sky130_fd_sc_hd__a22oi_1
XMuI._4695_ MuI._0209_ MuI._0261_ vssd1 vssd1 vccd1 vccd1 MuI._0408_ sky130_fd_sc_hd__xor2_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10499__A _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4906__A MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3646_ MuI._1307_ MuI._1802_ MuI._2440_ MuI._2451_ vssd1 vssd1 vccd1 vccd1 MuI._2462_
+ sky130_fd_sc_hd__and4_1
XMuI._6434_ MuI._2090_ MuI._2254_ MuI._2256_ MuI._2263_ vssd1 vssd1 vccd1 vccd1 MuI._2321_
+ sky130_fd_sc_hd__o31a_1
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09072__B _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _00237_ _00462_ _06431_ _00287_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__and4_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08133__A1 _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08133__B2 _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6365_ MuI._1930_ MuI._1936_ vssd1 vssd1 vccd1 vccd1 MuI._2245_ sky130_fd_sc_hd__or2b_1
XMuI._3577_ MuI._1648_ MuI._1692_ vssd1 vssd1 vccd1 vccd1 MuI._1703_ sky130_fd_sc_hd__and2_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08471_ _01074_ _01087_ _01083_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__nand3_1
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0955__B_N AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5316_ MuI._0959_ MuI._0957_ MuI._0958_ vssd1 vssd1 vccd1 vccd1 MuI._1091_ sky130_fd_sc_hd__or3_1
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4344__C MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6296_ MuI._2167_ MuI._2168_ vssd1 vssd1 vccd1 vccd1 MuI._2169_ sky130_fd_sc_hd__xor2_1
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _04703_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__buf_6
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3606__A1 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__B1 _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5247_ MuI._1009_ MuI._1011_ MuI._1013_ vssd1 vssd1 vccd1 vccd1 MuI._1015_ sky130_fd_sc_hd__and3_1
XANTENNA__07601__A _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07353_ _06652_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__nor2_1
XANTENNA__09633__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5178_ MuI._0937_ MuI._0938_ vssd1 vssd1 vccd1 vccd1 MuI._0939_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07320__B _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07284_ _02582_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4360__B MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4129_ MuI._3227_ MuI._3228_ vssd1 vssd1 vccd1 vccd1 MuI._3229_ sky130_fd_sc_hd__nand2_1
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _01638_ _01639_ _01633_ _01634_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a211o_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10962__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07947__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07947__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08789__D _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09925_ _02147_ _02159_ _02331_ _02332_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__o211a_1
XANTENNA__07048__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3704__B MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07990__B _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _02510_ _02501_ _02508_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__and3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06887__A _04208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08372__A1 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08372__B2 _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _02959_ _03960_ _06443_ _02905_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a22oi_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5295__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _02374_ _02435_ _02424_ _02434_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__o211a_1
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _05413_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[22\] sky130_fd_sc_hd__buf_2
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._3720__A MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _01354_ _01355_ _06680_ _00090_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__and4bb_1
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _01220_ _01286_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _06630_ _05380_ _06546_ _00012_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a22oi_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09710__B _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04473_ _04474_ _04250_ _04364_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__o211a_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _03343_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ _05724_ _02941_ _02731_ AuI.result\[27\] vssd1 vssd1 vccd1 vccd1 _06262_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5366__B MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _03243_ _03270_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__xnor2_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6011__A2 MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _02800_ _05141_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or2_1
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _06188_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nor2_1
X_10493_ _00727_ _04714_ _06613_ _00728_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__a22oi_1
XANTENNA__13184__A1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12232_ _05051_ _05067_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__or2_1
XFILLER_170_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08342__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A1 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11734__A2 _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1610_ AuI._0676_ AuI._0674_ vssd1 vssd1 vccd1 vccd1 AuI._0780_ sky130_fd_sc_hd__or2_1
X_12163_ _04864_ _04868_ _04993_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a211oi_1
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6197__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11114_ _03539_ _00678_ _00047_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__and3_1
XFILLER_150_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1541_ AuI._0652_ AuI._0657_ AuI._0658_ AuI._0647_ vssd1 vssd1 vccd1 vccd1 AuI._0723_
+ sky130_fd_sc_hd__a31o_1
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _04919_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__nor2_1
XFILLER_1_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11045_ _03606_ _03608_ _03607_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__o21bai_1
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1472_ AuI._0358_ AuI._0361_ vssd1 vssd1 vccd1 vccd1 AuI._0658_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06797__A _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6078__A2 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__B _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3500_ MuI._0812_ MuI._0845_ vssd1 vssd1 vccd1 vccd1 MuI._0856_ sky130_fd_sc_hd__xor2_2
XANTENNA__13239__A2 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4480_ MuI._2852_ MuI._2605_ MuI._3189_ MuI._2868_ vssd1 vssd1 vccd1 vccd1 MuI._0171_
+ sky130_fd_sc_hd__and4_1
XFILLER_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10112__A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _05887_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__xnor2_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3431_ MuI.a_operand\[30\] MuI.b_operand\[30\] vssd1 vssd1 vccd1 vccd1 MuI._0097_
+ sky130_fd_sc_hd__nand2_1
XFILLER_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _04761_ _04762_ _03133_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o21ai_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6150_ MuI._0328_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._2008_ sky130_fd_sc_hd__and2_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6786__B1 MuI._2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11878_ _04534_ _04536_ _04535_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__o21bai_1
XFILLER_177_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5101_ MuI._2765_ MuI._3402_ MuI._0020_ MuI._0477_ vssd1 vssd1 vccd1 vccd1 MuI._0854_
+ sky130_fd_sc_hd__a22oi_2
XMuI._6081_ MuI._1472_ MuI._1296_ MuI._1791_ MuI._2055_ vssd1 vssd1 vccd1 vccd1 MuI._1932_
+ sky130_fd_sc_hd__and4_1
XFILLER_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10829_ _03514_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__xor2_2
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5032_ MuI._0776_ MuI._0777_ vssd1 vssd1 vccd1 vccd1 MuI._0778_ sky130_fd_sc_hd__xor2_4
XFILLER_186_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4180__B MuI._3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1675__C1 AuI._0024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12981__B _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5707__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ _06391_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__or2_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__A1 _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5934_ MuI._1737_ MuI._1752_ vssd1 vssd1 vccd1 vccd1 MuI._1771_ sky130_fd_sc_hd__nor2_1
XANTENNA__07929__B2 _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._814_ AuI.pe._008_ AuI.pe._370_ AuI.pe._372_ AuI.pe._373_ AuI.pe._352_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._353_ sky130_fd_sc_hd__o41a_1
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5865_ MuI._1689_ MuI._1694_ vssd1 vssd1 vccd1 vccd1 MuI._1695_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07971_ _03335_ _04122_ _00300_ _00302_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3524__B1 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._745_ AuI.pe.significand\[21\] AuI.pe._270_ vssd1 vssd1 vccd1 vccd1 AuI.pe._290_
+ sky130_fd_sc_hd__nand2_1
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4816_ MuI._0536_ MuI._0538_ vssd1 vssd1 vccd1 vccd1 MuI._0541_ sky130_fd_sc_hd__or2b_1
X_09710_ _02377_ _06443_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__nand2_1
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06922_ _04585_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__buf_6
XMuI._5796_ MuI._1614_ MuI._1618_ vssd1 vssd1 vccd1 vccd1 MuI._1619_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._676_ AuI.pe._074_ AuI.pe._212_ AuI.pe._215_ AuI.pe._224_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[17\] sky130_fd_sc_hd__o22a_1
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4747_ MuI._0457_ MuI._0462_ MuI._0464_ vssd1 vssd1 vccd1 vccd1 MuI._0465_ sky130_fd_sc_hd__o21ai_1
X_09641_ _06520_ _06516_ net132 _06430_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and4_1
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06853_ _03842_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__and3_1
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13317__B _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4636__A MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12221__B _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3540__A MuI.b_operand\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4678_ MuI._0386_ MuI._0388_ vssd1 vssd1 vccd1 vccd1 MuI._0389_ sky130_fd_sc_hd__and2_1
XFuI._136__142 vssd1 vssd1 vccd1 vccd1 FuI._136__142/HI net142 sky130_fd_sc_hd__conb_1
X_09572_ _02177_ _02180_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06784_ _03099_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__buf_6
XMuI._6417_ MuI._2292_ MuI._2291_ vssd1 vssd1 vccd1 vccd1 MuI._2302_ sky130_fd_sc_hd__or2b_1
XFILLER_35_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3629_ MuI._2220_ MuI._2264_ vssd1 vssd1 vccd1 vccd1 MuI._2275_ sky130_fd_sc_hd__xor2_1
X_08523_ _00915_ _01140_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__nor2_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6348_ MuI._2224_ MuI._2225_ vssd1 vssd1 vccd1 vccd1 MuI._2226_ sky130_fd_sc_hd__nand2_1
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08454_ net119 _04294_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__nand2_1
XFILLER_211_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07405_ _00021_ _00022_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__nand2_1
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6279_ MuI._2057_ MuI._2060_ MuI._2058_ vssd1 vssd1 vccd1 vccd1 MuI._2150_ sky130_fd_sc_hd__o21ba_1
XFILLER_91_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4371__A MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ _00986_ _00987_ _01002_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__nand3_1
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07336_ _06617_ _06618_ _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21o_2
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4521__D MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07267_ _05241_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__buf_4
XFILLER_118_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _01437_ _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__and2_1
XFILLER_164_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07198_ _06475_ _05316_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nand2_1
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10206__A_N _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A2 _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09908_ _02524_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__xor2_1
XFILLER_120_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07506__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _06492_ _06463_ net127 _04100_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__and4_1
XFILLER_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09424__C _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07225__B _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__and2_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12781_ _05549_ _05601_ _05657_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__and3_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _04527_ _04528_ _04529_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o21ai_1
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4243__A1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11663_ _04454_ _04455_ _04457_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4243__B2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13402_ _06315_ _02915_ _02926_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__mux2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10614_ _03318_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._5096__B MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11594_ _04381_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
XFILLER_155_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11698__A _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A2 _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _06188_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__inv_2
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _03244_ _03252_ _03253_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__nand3_1
XFILLER_183_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0972_ net50 net18 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0184_ sky130_fd_sc_hd__mux2_1
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ _06171_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nor2_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10476_ _03140_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__xor2_2
XANTENNA__08072__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11210__B _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _05048_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__xnor2_1
XMuI._3980_ MuI._3075_ MuI._3076_ MuI._3079_ vssd1 vssd1 vccd1 vccd1 MuI._3080_ sky130_fd_sc_hd__a21bo_1
X_13195_ _05869_ _06039_ _03507_ _05992_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o211a_1
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._808__A AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6153__D1 MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ _04956_ _04975_ _04976_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__and3_1
XFILLER_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5262__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5650_ MuI._1290_ MuI._1457_ MuI._1288_ vssd1 vssd1 vccd1 vccd1 MuI._1458_ sky130_fd_sc_hd__o21ai_2
XAuI._1524_ AuI._0257_ AuI._0692_ vssd1 vssd1 vccd1 vccd1 AuI._0708_ sky130_fd_sc_hd__or2_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12077_ _04825_ _04827_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__or2_1
XAuI.pe._530_ AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 AuI.pe._089_ sky130_fd_sc_hd__clkbuf_4
XMuI._4601_ MuI.a_operand\[3\] vssd1 vssd1 vccd1 vccd1 MuI._0304_ sky130_fd_sc_hd__buf_2
XFILLER_38_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5581_ MuI._1379_ MuI._1380_ MuI._1381_ vssd1 vssd1 vccd1 vccd1 MuI._1382_ sky130_fd_sc_hd__o21a_1
X_11028_ _03771_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and3_1
XAuI._1455_ AuI._0451_ AuI._0454_ vssd1 vssd1 vccd1 vccd1 AuI._0641_ sky130_fd_sc_hd__and2b_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._461_ AuI.pe._025_ vssd1 vssd1 vccd1 vccd1 AuI.pe._026_ sky130_fd_sc_hd__buf_2
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4532_ MuI.a_operand\[4\] vssd1 vssd1 vccd1 vccd1 MuI._0228_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3809__B2 MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1386_ net18 net50 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0577_ sky130_fd_sc_hd__mux2_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._543__A AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4463_ MuI._0768_ MuI._3268_ MuI._0019_ MuI._0022_ vssd1 vssd1 vccd1 vccd1 MuI._0153_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12979_ _05868_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_1
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6202_ MuI._2028_ MuI._2064_ vssd1 vssd1 vccd1 vccd1 MuI._2065_ sky130_fd_sc_hd__xnor2_2
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4394_ MuI._0075_ MuI._0076_ vssd1 vssd1 vccd1 vccd1 MuI._0077_ sky130_fd_sc_hd__xor2_1
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10496__B _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6133_ MuI._1985_ MuI._1988_ vssd1 vssd1 vccd1 vccd1 MuI._1990_ sky130_fd_sc_hd__nor2_1
XFILLER_178_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6064_ MuI._1909_ MuI._1913_ vssd1 vssd1 vccd1 vccd1 MuI._1914_ sky130_fd_sc_hd__and2_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13396__B2 _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08170_ _00782_ _00787_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__xnor2_2
XANTENNA_MuI._3519__B MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5015_ MuI._0754_ MuI._0758_ MuI._0759_ MuI._0585_ vssd1 vssd1 vccd1 vccd1 MuI._0760_
+ sky130_fd_sc_hd__o211a_1
X_07121_ _06424_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4341__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1663__A2 AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07052_ _05981_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__buf_2
XFILLER_161_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 Exception sky130_fd_sc_hd__buf_2
XANTENNA__12216__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5917_ MuI._1740_ MuI._1751_ vssd1 vssd1 vccd1 vccd1 MuI._1752_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08710__A _00951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._6846__A MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5848_ MuI._2796_ MuI._3247_ MuI._0710_ MuI._0711_ vssd1 vssd1 vccd1 vccd1 MuI._1676_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07954_ _03002_ _00093_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__nand2_1
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._728_ AuI.pe._388_ AuI.pe._009_ vssd1 vssd1 vccd1 vccd1 AuI.pe._273_ sky130_fd_sc_hd__nand2_2
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4170__B1 MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06905_ _04391_ _04402_ _03766_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__and3_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5779_ MuI._0477_ MuI.a_operand\[10\] MuI._2866_ MuI._2868_ vssd1 vssd1 vccd1
+ vccd1 MuI._1600_ sky130_fd_sc_hd__and4_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07885_ _00502_ _03917_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__nand2_2
XANTENNA__11493__D _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11331__B1 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._659_ AuI.pe._372_ AuI.pe._141_ AuI.pe._201_ vssd1 vssd1 vccd1 vccd1 AuI.pe._209_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _02208_ _02257_ _02253_ _02256_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a211o_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06836_ _03658_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09541__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _02170_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a21o_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06767_ _02916_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__and3_1
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _00871_ _01122_ _01065_ _01120_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__o211a_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _06544_ _04358_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__nand2_1
XFILLER_196_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06698_ _02173_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[0\] sky130_fd_sc_hd__buf_2
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _01053_ _01052_ _01051_ _01007_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__o211a_1
XFILLER_197_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._141_ FuI._003_ net147 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[12\] sky130_fd_sc_hd__dlxtn_1
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11014__C _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ _00970_ _00984_ _00985_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__nand3_2
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._072_ FuI._036_ FuI._037_ FuI._038_ FuI._039_ FuI._035_ vssd1 vssd1 vccd1 vccd1
+ FuI._040_ sky130_fd_sc_hd__a41o_1
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ net39 vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__buf_6
XFILLER_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08299_ _00605_ _00604_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__and2b_1
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08604__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ _01147_ _01146_ _04649_ _04714_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__and4_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12126__B _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ AuI.result\[1\] _02938_ _02940_ _02942_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12000_ _03658_ _00550_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nand2_1
XANTENNA__09716__A _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _02826_ _02842_ _02857_ _02872_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__or4b_1
XFILLER_79_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09435__B _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07236__A net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0917__A1 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _00290_ _00289_ _03247_ _00783_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__and4_1
XAuI._1240_ AuI._0420_ AuI._0442_ vssd1 vssd1 vccd1 vccd1 AuI._0443_ sky130_fd_sc_hd__nand2_1
XANTENNA__11873__A1 _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__B2 _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _03733_ _05327_ _05637_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nand3_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1171_ net32 net64 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0378_ sky130_fd_sc_hd__mux2_2
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09818__A1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05517_ _05518_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and2_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08067__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6205__A2 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _04374_ _04377_ _04375_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o21bai_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _05565_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._5538__C MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11646_ _03722_ _04660_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and2_2
XFILLER_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 a_operand[18] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_6
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput25 a_operand[28] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_4
Xinput36 a_operand[9] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
X_11577_ _04250_ _04252_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nand4_2
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 b_operand[19] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10061__B1 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput58 b_operand[29] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_4
X_13316_ _03561_ _03626_ _05906_ _05981_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and4_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10528_ _03231_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__a21o_1
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0955_ AuI._0166_ AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 AuI._0167_ sky130_fd_sc_hd__or2b_1
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6820_ MuI._2707_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2741_ sky130_fd_sc_hd__and2_1
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13247_ _06151_ _06152_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__o21a_1
XFILLER_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ _02984_ _04520_ _00036_ _02983_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__a22o_1
XAuI._0886_ AuI._0096_ AuI._0097_ AuI._0099_ AuI._0105_ vssd1 vssd1 vccd1 vccd1 AuI._0106_
+ sky130_fd_sc_hd__and4bb_1
XMuI._6751_ MuI._2505_ MuI._2664_ vssd1 vssd1 vccd1 vccd1 MuI._2669_ sky130_fd_sc_hd__nand2_1
XMuI._3963_ MuI._2981_ MuI._2988_ vssd1 vssd1 vccd1 vccd1 MuI._3063_ sky130_fd_sc_hd__nand2_1
X_13178_ _03400_ _05531_ _02743_ _02736_ MuI.result\[24\] vssd1 vssd1 vccd1 vccd1
+ _06085_ sky130_fd_sc_hd__a32o_1
XFILLER_123_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11875__B _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5702_ MuI._1512_ MuI._1513_ MuI._1514_ vssd1 vssd1 vccd1 vccd1 MuI._1515_ sky130_fd_sc_hd__or3_1
XFILLER_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6682_ MuI._0013_ MuI._2592_ vssd1 vssd1 vccd1 vccd1 MuI._2593_ sky130_fd_sc_hd__xnor2_1
X_12129_ _04792_ _04801_ _04799_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__o21bai_1
XMuI._3894_ MuI._2990_ MuI._2991_ MuI._2992_ MuI._2993_ vssd1 vssd1 vccd1 vccd1 MuI._2994_
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A1 _00918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5633_ MuI._3269_ MuI._0421_ MuI._1415_ MuI._1416_ vssd1 vssd1 vccd1 vccd1 MuI._1440_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13302__A1 _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1507_ AuI._0692_ vssd1 vssd1 vccd1 vccd1 AuI._0693_ sky130_fd_sc_hd__buf_2
XANTENNA__07146__A _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._513_ AuI.pe._072_ AuI.pe._065_ vssd1 vssd1 vccd1 vccd1 AuI.pe._073_ sky130_fd_sc_hd__nand2_1
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5564_ MuI._1361_ MuI._1363_ vssd1 vssd1 vccd1 vccd1 MuI._1364_ sky130_fd_sc_hd__nor2_1
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1030__A0 net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1438_ AuI._0473_ AuI._0477_ vssd1 vssd1 vccd1 vccd1 AuI._0624_ sky130_fd_sc_hd__and2_1
XANTENNA__10667__A2 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _00278_ _03432_ _06431_ _00287_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__and4_1
XANTENNA__06985__A _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._444_ AuI.pe.significand\[5\] AuI.pe._010_ vssd1 vssd1 vccd1 vccd1 AuI.pe._011_
+ sky130_fd_sc_hd__and2b_1
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4515_ MuI.b_operand\[14\] MuI._2352_ vssd1 vssd1 vccd1 vccd1 MuI._0210_ sky130_fd_sc_hd__nand2_1
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5495_ MuI._1183_ MuI._1242_ MuI._1287_ vssd1 vssd1 vccd1 vccd1 MuI._1288_ sky130_fd_sc_hd__or3_1
XFILLER_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1369_ AuI._0257_ AuI._0558_ AuI._0559_ AuI._0560_ vssd1 vssd1 vccd1 vccd1 AuI._0562_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09809__A1 _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__B2 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4446_ MuI._0132_ MuI._0133_ vssd1 vssd1 vccd1 vccd1 MuI._0134_ sky130_fd_sc_hd__xor2_1
X_09340_ _01924_ _01956_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09080__B _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4377_ MuI._0056_ MuI._0058_ vssd1 vssd1 vccd1 vccd1 MuI._0059_ sky130_fd_sc_hd__or2b_1
XFILLER_178_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _01779_ _01884_ _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._5404__B1 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6116_ MuI._1021_ MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 MuI._1971_ sky130_fd_sc_hd__nand2_2
XANTENNA__11830__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08222_ _06560_ _04972_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__nand2_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10954__B _03655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6047_ MuI._0779_ MuI._1021_ MuI._2704_ MuI._2649_ vssd1 vssd1 vccd1 vccd1 MuI._1895_
+ sky130_fd_sc_hd__and4_1
XANTENNA_AuI._1356__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _00399_ _00400_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout122_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07104_ _05338_ _06414_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__and2_1
XFILLER_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08084_ _00700_ _00698_ _00699_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__nand3_2
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07035_ _05799_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[28\] sky130_fd_sc_hd__clkbuf_2
XFILLER_106_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._448__A AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07220__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08986_ _01467_ _01461_ _01466_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a21o_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07937_ _00011_ _06612_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__and2_4
XANTENNA_MuI._3497__A2 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11855__A1 _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07868_ _00270_ _04369_ _00232_ _00230_ _04456_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a32o_1
XANTENNA__11855__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09607_ _02199_ _02197_ _02198_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__or3_1
X_06819_ net55 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__buf_4
XFILLER_84_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07799_ _00413_ _00415_ _00411_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11306__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09538_ _02604_ _02669_ _03873_ _03971_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__and4_1
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09276__A2 _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _02205_ _00035_ _00030_ _06534_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a22oi_2
XFILLER_106_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ _04280_ _04278_ _04279_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__nand3_2
XFILLER_169_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4749__A2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _05333_ _05334_ _05226_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__o21ai_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFuI._124_ FuI._061_ FuI._026_ net105 FuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1
+ FuI._009_ sky130_fd_sc_hd__o211a_1
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08615__A _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3957__B1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _04075_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__nor3_1
XANTENNA_AuI._1088__A0 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08236__B1 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11041__A _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12583__A2 _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _04113_ _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nand3_1
XFILLER_192_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10594__A1 _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10594__B2 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _02782_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._6189__C MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10313_ _02957_ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__xor2_2
XANTENNA__11976__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ _00058_ _05391_ _04056_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__a22o_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13032_ _02779_ _05927_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or2_1
XANTENNA_input52_A b_operand[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10244_ _02755_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__xnor2_1
XFILLER_106_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09446__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6659__C1 MuI._2563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12797__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09165__B _01722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10175_ _03067_ _05134_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__or2_1
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12099__A1 _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12099__B2 _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5540__D MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1012__A0 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1223_ AuI._0420_ AuI._0425_ AuI._0426_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0427_
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4300_ MuI._3263_ MuI._3398_ vssd1 vssd1 vccd1 vccd1 MuI._3400_ sky130_fd_sc_hd__and2_1
XMuI._5280_ MuI._1048_ MuI._1049_ MuI._1029_ vssd1 vssd1 vccd1 vccd1 MuI._1051_ sky130_fd_sc_hd__a21oi_2
XAuI._1154_ AuI._0256_ AuI._0359_ AuI._0360_ AuI._0361_ vssd1 vssd1 vccd1 vccd1 AuI._0362_
+ sky130_fd_sc_hd__and4_1
X_12816_ _05617_ _05619_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__nand2_1
XANTENNA__07413__B _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09267__A2 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4231_ MuI._3198_ MuI._3330_ vssd1 vssd1 vccd1 vccd1 MuI._3331_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _05614_ _05620_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nand3_1
XAuI._1085_ AuI._0153_ AuI._0295_ AuI._0212_ vssd1 vssd1 vccd1 vccd1 AuI._0296_ sky130_fd_sc_hd__a21o_1
XFILLER_188_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4162_ MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 MuI._3262_ sky130_fd_sc_hd__buf_4
XFILLER_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12678_ _05419_ _05547_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or3_1
XFILLER_175_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4093_ MuI._3191_ MuI._3192_ vssd1 vssd1 vccd1 vccd1 MuI._3193_ sky130_fd_sc_hd__nor2_1
X_11629_ _04418_ _04419_ _04385_ _04244_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__a211oi_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12047__A _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10585__A1 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0938_ AuI._0147_ AuI._0149_ AuI._0097_ vssd1 vssd1 vccd1 vccd1 AuI._0150_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI.pe._558__A2 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6803_ MuI._2695_ MuI._2717_ MuI._2718_ MuI._2725_ vssd1 vssd1 vccd1 vccd1 MuI._2727_
+ sky130_fd_sc_hd__and4_1
XFILLER_171_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08898__C _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4995_ MuI._0643_ MuI._0639_ vssd1 vssd1 vccd1 vccd1 MuI._0738_ sky130_fd_sc_hd__and2b_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08260__A _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0869_ AuI._0072_ AuI._0073_ AuI._0069_ vssd1 vssd1 vccd1 vccd1 AuI._0089_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6734_ MuI._2444_ MuI._2648_ MuI._2468_ vssd1 vssd1 vccd1 vccd1 MuI._2651_ sky130_fd_sc_hd__o21a_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6114__A1 MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3946_ MuI._3043_ MuI._3044_ MuI._3045_ vssd1 vssd1 vccd1 vccd1 MuI._3046_ sky130_fd_sc_hd__nand3_1
X_08840_ _06463_ net133 _06581_ _02107_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a22o_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4125__B1 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6665_ MuI._2570_ MuI._2574_ MuI._2485_ vssd1 vssd1 vccd1 vccd1 MuI._2575_ sky130_fd_sc_hd__mux2_1
XFILLER_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3877_ MuI._1010_ MuI._2975_ MuI._2976_ MuI._0779_ vssd1 vssd1 vccd1 vccd1 MuI._2977_
+ sky130_fd_sc_hd__a22oi_2
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _02948_ _06430_ _06431_ _00028_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__a22o_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5616_ MuI._1415_ MuI._1418_ MuI._1420_ vssd1 vssd1 vccd1 vccd1 MuI._1421_ sky130_fd_sc_hd__o21a_1
X_07722_ _00069_ _00106_ _00144_ _00145_ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a211oi_1
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6596_ MuI._0196_ MuI._0185_ MuI._0163_ vssd1 vssd1 vccd1 vccd1 MuI._2499_ sky130_fd_sc_hd__and3b_1
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11837__B2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5547_ MuI._1311_ MuI._1310_ MuI._1302_ vssd1 vssd1 vccd1 vccd1 MuI._1345_ sky130_fd_sc_hd__a21o_1
XFILLER_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07653_ net125 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkbuf_4
XAuI.pe._427_ AuI.pe.significand\[9\] AuI.pe.significand\[10\] AuI.pe.significand\[11\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._394_ sky130_fd_sc_hd__nor3_1
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11126__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5478_ MuI._1260_ MuI._1267_ MuI._1268_ vssd1 vssd1 vccd1 vccd1 MuI._1269_ sky130_fd_sc_hd__nand3_1
XANTENNA__07323__B _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5459__B MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07584_ _00195_ _00196_ _00201_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__nand3_1
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4429_ MuI._0105_ MuI._0114_ vssd1 vssd1 vccd1 vccd1 MuI._0115_ sky130_fd_sc_hd__and2_1
X_09323_ _01940_ _01894_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09254_ _01653_ _01869_ _01870_ _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_167_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10684__B _06605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ _06475_ _06525_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5475__A MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__A1 _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09185_ _02808_ _06443_ _00303_ _02765_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12014__B2 _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ _02840_ _00423_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5194__B MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ _06429_ _04057_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3426__C MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07018_ net23 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11525__B1 _04308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12813__A1_N _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4667__A1 MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4667__B2 MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _01585_ _01584_ _01530_ _01528_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__o211ai_2
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11828__A1 _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ _04684_ _04686_ _04685_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__o21bai_1
XANTENNA__12420__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _02544_ _02554_ _02563_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07514__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09432__C _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _03393_ _03413_ _03591_ _03592_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a211oi_4
XFILLER_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4273__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ _05422_ _05326_ _05464_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__o211a_1
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3642__A2 MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10875__A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _06442_ _00093_ _04520_ _06444_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a22oi_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ MuI.result\[17\] _02738_ _02931_ FuI.Integer\[17\] _05390_ vssd1 vssd1 vccd1
+ vccd1 _05392_ sky130_fd_sc_hd__a221o_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6041__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ _05311_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__xor2_1
XFILLER_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13202__B1 _05906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._107_ FuI._052_ FuI._060_ FuI._063_ FuI.a_operand\[12\] vssd1 vssd1 vccd1 vccd1
+ FuI._002_ sky130_fd_sc_hd__o31a_1
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _00216_ _03051_ _05574_ _00217_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__a22o_1
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _05240_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI._0808__B1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _03966_ _03977_ _03976_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__a21o_1
XANTENNA__07432__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07432__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11276_ _03927_ _03930_ _03929_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__o21bai_1
XFILLER_140_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3800_ MuI._2894_ MuI._0768_ MuI._2867_ MuI._2869_ vssd1 vssd1 vccd1 vccd1 MuI._2900_
+ sky130_fd_sc_hd__and4_1
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11856__D _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _05908_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and2_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4780_ MuI._0312_ MuI._0498_ MuI._0497_ vssd1 vssd1 vccd1 vccd1 MuI._0501_ sky130_fd_sc_hd__o21a_1
XANTENNA__09185__B2 _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ _03507_ _05671_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__and2b_1
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3731_ MuI._2830_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._2831_ sky130_fd_sc_hd__nand2_1
XANTENNA_AuI.pe._816__A AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10158_ _03454_ _05595_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__and2b_1
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6450_ MuI._2331_ MuI._2336_ MuI._2309_ vssd1 vssd1 vccd1 vccd1 MuI._2338_ sky130_fd_sc_hd__o21a_1
XMuI._3662_ MuI.b_operand\[12\] vssd1 vssd1 vccd1 vccd1 MuI._2638_ sky130_fd_sc_hd__buf_2
XFILLER_208_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10089_ _04186_ _02345_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__and2b_1
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5401_ MuI._1137_ MuI._1128_ MuI._1136_ vssd1 vssd1 vccd1 vccd1 MuI._1184_ sky130_fd_sc_hd__nand3_1
XANTENNA__10769__B _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6381_ MuI._2260_ MuI._2261_ vssd1 vssd1 vccd1 vccd1 MuI._2262_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3593_ MuI._1340_ MuI._1868_ vssd1 vssd1 vccd1 vccd1 MuI._1879_ sky130_fd_sc_hd__nor2_1
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5332_ MuI._1107_ vssd1 vssd1 vccd1 vccd1 MuI._1108_ sky130_fd_sc_hd__inv_2
XFILLER_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1206_ AuI._0407_ AuI._0409_ AuI._0410_ AuI._0288_ AuI._0249_ vssd1 vssd1 vccd1
+ vccd1 AuI._0411_ sky130_fd_sc_hd__a221o_2
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4183__B MuI._3171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5263_ MuI._2484_ MuI._2885_ MuI._2881_ MuI._0327_ vssd1 vssd1 vccd1 vccd1 MuI._1033_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1137_ net30 net62 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0346_ sky130_fd_sc_hd__mux2_1
XFILLER_188_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4214_ MuI._3313_ MuI._3193_ vssd1 vssd1 vccd1 vccd1 MuI._3314_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5194_ MuI._3349_ MuI._3268_ vssd1 vssd1 vccd1 vccd1 MuI._0957_ sky130_fd_sc_hd__nand2_1
XFILLER_176_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1068_ AuI._0237_ AuI._0278_ AuI._0175_ vssd1 vssd1 vccd1 vccd1 AuI._0279_ sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__C _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4145_ MuI.a_operand\[4\] vssd1 vssd1 vccd1 vccd1 MuI._3245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3808__A MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4076_ MuI._3158_ MuI._3175_ vssd1 vssd1 vccd1 vccd1 MuI._3176_ sky130_fd_sc_hd__xor2_1
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5543__C1 MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09086__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5742__B MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ _02598_ _02600_ _02601_ _02602_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a211o_1
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12704__C1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3543__A MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1224__A0 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4978_ MuI._1274_ MuI._0245_ MuI._0717_ MuI._0718_ vssd1 vssd1 vccd1 vccd1 MuI._0719_
+ sky130_fd_sc_hd__a31o_1
X_09872_ _02527_ _02512_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__or2_1
XFILLER_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4358__B MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6717_ MuI._2588_ MuI._2597_ MuI._2601_ MuI._2631_ vssd1 vssd1 vccd1 vccd1 MuI._2632_
+ sky130_fd_sc_hd__and4_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07726__A2 _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3929_ MuI._2935_ MuI._2936_ vssd1 vssd1 vccd1 vccd1 MuI._3029_ sky130_fd_sc_hd__or2_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08823_ _01438_ _01439_ _01440_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__or3_1
XFILLER_86_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__A1 _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__B2 _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6648_ MuI._3403_ MuI._0421_ MuI._1414_ MuI._1441_ vssd1 vssd1 vccd1 vccd1 MuI._2556_
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _01369_ _01371_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__and2b_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07334__A _06629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07705_ _03432_ _04165_ _04229_ net113 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__a22o_1
XMuI._6579_ MuI._2478_ MuI._0988_ MuI._0394_ MuI._0548_ vssd1 vssd1 vccd1 vccd1 MuI._2480_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _01017_ _01018_ _01048_ _01049_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__or4bb_2
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _00252_ _00212_ _00213_ _00251_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__and4_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5074__A1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5074__B2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07567_ _00171_ _00172_ _00183_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__and3_2
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09306_ _01913_ _01915_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10246__B1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07498_ _03013_ _04660_ _00065_ _00061_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__a31o_1
XANTENNA__08165__A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _01631_ _01852_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__o211a_1
XFILLER_210_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4585__B1 MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09168_ _06579_ _00266_ _00592_ _02582_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5355__D MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _00734_ _00735_ _00736_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__or3_1
X_09099_ _01714_ _01715_ _01716_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__or3_1
XFILLER_107_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11957__C _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11130_ _03757_ _03760_ _03758_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21bai_1
XANTENNA_MuI._4549__A MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__C net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09167__A1 _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__B _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3453__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _03632_ _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__xor2_1
XFILLER_89_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ _01202_ _01318_ _01317_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a21oi_1
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10721__A1 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__B2 _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09879__A1_N _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13246__A _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A a_operand[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07244__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3863__A2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11963_ _04665_ _04667_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__nand2_1
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4715__C MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ _03647_ _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__xnor2_2
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ _03744_ _04725_ _04563_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nand3_1
XFILLER_205_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10845_ _03574_ _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nor2_1
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6703__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10776_ _02750_ _03327_ _03487_ _03488_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__a221o_1
XFILLER_185_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10788__A1 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4731__B MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__B1 _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12515_ _05363_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__nor2_1
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11213__B _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13495_ _02812_ _02820_ _06365_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__or3_1
XFILLER_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__A2 _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ _03722_ _05123_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nand2_1
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5950_ MuI._1782_ MuI._1786_ MuI._1787_ vssd1 vssd1 vccd1 vccd1 MuI._1788_ sky130_fd_sc_hd__nand3b_1
XFILLER_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _05180_ _05224_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__or3_2
XAuI.pe._830_ AuI.operand_a\[29\] AuI.pe._365_ vssd1 vssd1 vccd1 vccd1 AuI.exponent_sub\[6\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4901_ MuI._0631_ MuI._0621_ MuI._0629_ vssd1 vssd1 vccd1 vccd1 MuI._0634_ sky130_fd_sc_hd__nand3_1
XFILLER_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5881_ MuI._1646_ MuI._1711_ vssd1 vssd1 vccd1 vccd1 MuI._1712_ sky130_fd_sc_hd__xnor2_1
XANTENNA_output83_A net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _03898_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__inv_2
XFILLER_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._761_ AuI.pe._385_ AuI.pe.significand\[20\] AuI.pe._384_ AuI.pe._386_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._305_ sky130_fd_sc_hd__o211a_1
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12044__B _04866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4832_ MuI._0506_ MuI._0557_ vssd1 vssd1 vccd1 vccd1 MuI._0558_ sky130_fd_sc_hd__nor2_1
XFILLER_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11259_ _02566_ _03315_ _03849_ _04022_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__a31o_2
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._692_ AuI.pe._238_ AuI.pe._239_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._240_
+ sky130_fd_sc_hd__a21o_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08905__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4763_ MuI._2841_ MuI._2773_ MuI._0329_ MuI._0330_ vssd1 vssd1 vccd1 vccd1 MuI._0483_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08905__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6502_ MuI._2384_ MuI._2394_ vssd1 vssd1 vccd1 vccd1 MuI._2395_ sky130_fd_sc_hd__or2b_1
XMuI._3714_ MuI.b_operand\[19\] vssd1 vssd1 vccd1 vccd1 MuI._2814_ sky130_fd_sc_hd__buf_2
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4694_ MuI._0403_ MuI._0404_ MuI._0406_ vssd1 vssd1 vccd1 vccd1 MuI._0407_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6433_ MuI._2282_ MuI._2310_ MuI._2318_ vssd1 vssd1 vccd1 vccd1 MuI._2320_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._4906__B MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._697__A1 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__B _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3645_ MuI.a_operand\[12\] vssd1 vssd1 vccd1 vccd1 MuI._2451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09072__C net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12995__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6364_ MuI._2102_ MuI._2103_ MuI._2106_ vssd1 vssd1 vccd1 vccd1 MuI._2244_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4625__C MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08133__A2 _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3576_ MuI._1593_ MuI._1615_ MuI._1637_ vssd1 vssd1 vccd1 vccd1 MuI._1692_ sky130_fd_sc_hd__a21o_1
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _01074_ _01083_ _01087_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__a21o_1
XFILLER_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6253__B1 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5315_ MuI._1088_ MuI._1089_ vssd1 vssd1 vccd1 vccd1 MuI._1090_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07421_ _06599_ _06611_ _04832_ _06598_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a22o_1
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4344__D MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6295_ MuI._2131_ MuI._2104_ MuI._2135_ vssd1 vssd1 vccd1 vccd1 MuI._2168_ sky130_fd_sc_hd__a21oi_2
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12217__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3606__A2 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12217__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5246_ MuI._1009_ MuI._1011_ MuI._1013_ vssd1 vssd1 vccd1 vccd1 MuI._1014_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07601__B _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07352_ _06500_ _05563_ _05638_ _06501_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__a22oi_1
XFILLER_204_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__A2 _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3538__A MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5177_ MuI._0815_ MuI._0817_ MuI._0816_ vssd1 vssd1 vccd1 vccd1 MuI._0938_ sky130_fd_sc_hd__o21ba_1
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07283_ _06581_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__buf_4
XFILLER_176_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A_N _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4360__C MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4128_ MuI._3219_ MuI._3221_ vssd1 vssd1 vccd1 vccd1 MuI._3228_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _01633_ _01634_ _01638_ _01639_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__o211ai_2
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11728__B1 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10962__B _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4059_ MuI._2994_ MuI._3077_ MuI._3078_ vssd1 vssd1 vccd1 vccd1 MuI._3159_ sky130_fd_sc_hd__o21ai_1
XFILLER_191_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07947__A2 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__A _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09924_ _01959_ _01964_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__or2b_1
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3704__C MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input7_A a_operand[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _02501_ _02508_ _02510_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a21o_1
XFILLER_112_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07990__C _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13066__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08372__A2 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08806_ _00049_ _00062_ _06436_ _04035_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__and4_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5295__A1 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06998_ _05402_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__and3_1
X_09786_ _02424_ _02434_ _02374_ _02435_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a211oi_2
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5295__B2 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07064__A _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3720__B MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11259__A2 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _06622_ _04434_ _00098_ _00414_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__a22oi_1
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10202__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _01221_ _01222_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__nor2_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12504__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ net118 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__clkbuf_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _01215_ _01216_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__nor2_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ _02965_ _04316_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__nand2_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09085__B1 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3448__A MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ _03266_ _03269_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__xor2_2
XFILLER_195_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08832__B1 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _02800_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nand2_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _06189_ _06187_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__nor2_1
XFILLER_155_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10492_ _03192_ _03193_ _03194_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21o_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ _05051_ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nand2_1
XFILLER_170_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08342__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07938__A2 _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12162_ _04991_ _04992_ _04902_ _04903_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__o211a_1
XFILLER_163_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _03713_ _03731_ _03732_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__and3_1
XANTENNA__08061__C _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1540_ AuI._0606_ AuI._0720_ AuI._0722_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[3\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12093_ _03228_ _03282_ _05445_ _05509_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__and4_1
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4730__B1 MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _03786_ _03787_ _03788_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__o21ai_1
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1471_ AuI._0653_ AuI._0654_ AuI._0655_ AuI._0656_ vssd1 vssd1 vccd1 vccd1 AuI._0657_
+ sky130_fd_sc_hd__a211o_1
XFILLER_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1303__A AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09173__B _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12995_ _03669_ _05585_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nand2_1
XMuI._3430_ MuI.a_operand\[30\] MuI.b_operand\[30\] vssd1 vssd1 vccd1 vccd1 MuI._0086_
+ sky130_fd_sc_hd__or2_2
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11946_ _04612_ _04613_ _04620_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o21ba_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5100_ MuI._2785_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0853_ sky130_fd_sc_hd__nand2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _04684_ _04685_ _04686_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6080_ MuI._2473_ MuI._3091_ vssd1 vssd1 vccd1 vccd1 MuI._1931_ sky130_fd_sc_hd__nand2_1
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ _03516_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4461__B MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5031_ MuI._0656_ MuI._0662_ vssd1 vssd1 vccd1 vccd1 MuI._0777_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11958__B1 _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10759_ _03479_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__xnor2_4
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _01330_ _06374_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12429_ _05164_ _05167_ _05165_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o21bai_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5933_ MuI._1731_ MuI._1733_ vssd1 vssd1 vccd1 vccd1 MuI._1770_ sky130_fd_sc_hd__nand2_1
XANTENNA__07929__A2 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07149__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._813_ AuI.pe._368_ AuI.pe._369_ AuI.pe._347_ AuI.pe._351_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._352_ sky130_fd_sc_hd__or4_1
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5864_ MuI._1690_ MuI._1693_ vssd1 vssd1 vccd1 vccd1 MuI._1694_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11894__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _00564_ _00586_ _00587_ _00339_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__o211a_1
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3524__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._744_ AuI.pe._059_ AuI.pe._213_ AuI.pe._284_ AuI.pe._288_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._289_ sky130_fd_sc_hd__a211o_1
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06988__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4815_ MuI._0422_ MuI._0500_ vssd1 vssd1 vccd1 vccd1 MuI._0540_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._3524__B2 MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ _04574_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__buf_4
XMuI._5795_ MuI._1616_ MuI._1617_ vssd1 vssd1 vccd1 vccd1 MuI._1618_ sky130_fd_sc_hd__nor2_1
XFILLER_141_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1669_ AuI._0702_ AuI._0697_ vssd1 vssd1 vccd1 vccd1 AuI._0021_ sky130_fd_sc_hd__or2_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._675_ AuI.pe._106_ AuI.pe._097_ AuI.pe._217_ AuI.pe._219_ AuI.pe._223_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._224_ sky130_fd_sc_hd__a2111o_1
XFILLER_110_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4746_ MuI._0351_ MuI._0463_ vssd1 vssd1 vccd1 vccd1 MuI._0464_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09640_ _02229_ _06436_ _06446_ _02431_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22oi_1
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06852_ _03831_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__buf_4
XANTENNA__10158__A_N _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__A _02991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4636__B MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4677_ MuI._0346_ MuI._0387_ vssd1 vssd1 vccd1 vccd1 MuI._0388_ sky130_fd_sc_hd__nor2_1
X_09571_ _02189_ _02190_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nand3_2
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06783_ net117 vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__buf_4
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6416_ MuI._2299_ MuI._2296_ vssd1 vssd1 vccd1 vccd1 MuI._2301_ sky130_fd_sc_hd__xor2_1
XMuI._3628_ MuI._2231_ MuI._2253_ vssd1 vssd1 vccd1 vccd1 MuI._2264_ sky130_fd_sc_hd__and2_1
X_08522_ _00914_ _00911_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__and2b_1
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6347_ MuI._2217_ MuI._2223_ vssd1 vssd1 vccd1 vccd1 MuI._2225_ sky130_fd_sc_hd__or2_1
XANTENNA__07612__A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5748__A MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3559_ MuI._1494_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._1505_ sky130_fd_sc_hd__nand2_1
X_08453_ net120 net44 _00089_ _00082_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__and4_1
XFILLER_23_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07404_ _00020_ _00019_ _06679_ _06678_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__a211o_1
XANTENNA__11134__A _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6278_ MuI._2146_ MuI._2148_ vssd1 vssd1 vccd1 vccd1 MuI._2149_ sky130_fd_sc_hd__xor2_1
XFILLER_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _00992_ _01001_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__xor2_1
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5229_ MuI._2841_ MuI._0228_ vssd1 vssd1 vccd1 vccd1 MuI._0995_ sky130_fd_sc_hd__nand2_1
XFILLER_177_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07335_ _06628_ _06635_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1428__B_N AuI._0550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _06560_ _06561_ _06563_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__nand4_1
X_09005_ _01410_ _01415_ _01436_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__or3_1
XFILLER_118_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07197_ _06486_ _06487_ _06497_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a21o_1
XFILLER_117_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07059__A _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5504__A2 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06898__A _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09907_ _02516_ _02545_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or2b_1
XFILLER_120_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3731__A MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A1 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11309__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _02477_ _02478_ _02469_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__a21o_1
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09424__D _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _00150_ net125 _00266_ _06469_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a22oi_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4265__C MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _04602_ _04603_ _04475_ _04497_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a211o_1
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__C _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12780_ _05549_ _05601_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__a21oi_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11731_ _04527_ _04528_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__or3_1
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _04275_ _04277_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__nand2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ _02829_ _06218_ _02828_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o21ba_1
X_10613_ _03323_ _03325_ _02926_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__mux2_1
XFILLER_211_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5096__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11593_ _04230_ _04366_ _04379_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__nor3_1
XFILLER_183_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1657__B1 AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ _03249_ _03251_ _03245_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a21o_1
X_13332_ _06241_ _06242_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__or2_1
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0971_ AuI._0180_ AuI._0182_ AuI._0176_ vssd1 vssd1 vccd1 vccd1 AuI._0183_ sky130_fd_sc_hd__mux2_1
XFILLER_182_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10475_ _03157_ _03177_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__xnor2_2
X_13263_ _06170_ _06168_ _06169_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__and3b_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08072__B _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12214_ _04913_ _04914_ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13194_ _06052_ _06050_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6153__C1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _04973_ _04974_ _04957_ _04847_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211ai_1
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1523_ AuI._0606_ AuI._0706_ AuI._0707_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[1\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09184__A _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5840__B MuI._1666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _02848_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4600_ MuI.b_operand\[19\] MuI.b_operand\[18\] MuI._0228_ MuI._3371_ vssd1 vssd1
+ vccd1 vccd1 MuI._0303_ sky130_fd_sc_hd__and4_1
XFILLER_110_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5580_ MuI._2882_ MuI._0315_ MuI._0320_ MuI._2886_ vssd1 vssd1 vccd1 vccd1 MuI._1381_
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ _03754_ _03756_ _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21oi_2
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1454_ AuI._0635_ AuI._0636_ AuI._0637_ AuI._0638_ AuI._0639_ vssd1 vssd1 vccd1
+ vccd1 AuI._0640_ sky130_fd_sc_hd__o2111a_1
XAuI.pe._460_ AuI.pe.significand\[23\] vssd1 vssd1 vccd1 vccd1 AuI.pe._025_ sky130_fd_sc_hd__buf_2
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4531_ MuI._0215_ MuI._0223_ MuI._0225_ vssd1 vssd1 vccd1 vccd1 MuI._0227_ sky130_fd_sc_hd__and3_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3809__A2 MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1385_ AuI._0375_ AuI._0498_ AuI._0574_ vssd1 vssd1 vccd1 vccd1 AuI._0576_ sky130_fd_sc_hd__o21ai_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4462_ MuI._1021_ MuI._3269_ MuI._0149_ MuI._0150_ vssd1 vssd1 vccd1 vccd1 MuI._0151_
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._521__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6201_ MuI._2030_ MuI._2029_ vssd1 vssd1 vccd1 vccd1 MuI._2064_ sky130_fd_sc_hd__nor2_1
X_12978_ _03389_ _05831_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__and3_1
XANTENNA__08528__A _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4393_ MuI._3392_ MuI._3416_ vssd1 vssd1 vccd1 vccd1 MuI._0076_ sky130_fd_sc_hd__xnor2_2
XFILLER_206_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11929_ _04547_ _04549_ _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__o211a_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6132_ MuI._1986_ MuI._1987_ vssd1 vssd1 vccd1 vccd1 MuI._1988_ sky130_fd_sc_hd__and2_1
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6063_ MuI._3154_ MuI._1842_ MuI._1908_ vssd1 vssd1 vccd1 vccd1 MuI._1913_ sky130_fd_sc_hd__or3_1
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13396__A2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3519__C MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1648__B1 AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5014_ MuI._0572_ MuI._0573_ MuI._0584_ vssd1 vssd1 vccd1 vccd1 MuI._0759_ sky130_fd_sc_hd__a21o_1
X_07120_ _05853_ _06414_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__and2_1
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5195__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3816__A MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ _05970_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 Overflow sky130_fd_sc_hd__buf_2
XFILLER_115_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__B1 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5916_ MuI._1749_ MuI._1750_ vssd1 vssd1 vccd1 vccd1 MuI._1751_ sky130_fd_sc_hd__or2b_1
XFILLER_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__B_N _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__A _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__B _00953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5847_ MuI._1673_ MuI._1674_ vssd1 vssd1 vccd1 vccd1 MuI._1675_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._6846__B MuI._2733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07973__A2_N _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _02894_ _02948_ _00098_ _00047_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__and4_1
XAuI.pe._727_ AuI.pe._258_ AuI.pe._269_ AuI.pe._272_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[20\]
+ sky130_fd_sc_hd__o21a_1
XMuI._5778_ MuI._0168_ MuI._3223_ vssd1 vssd1 vccd1 vccd1 MuI._1599_ sky130_fd_sc_hd__nand2_1
X_06904_ _02031_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__clkbuf_2
X_07884_ net61 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11331__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._658_ AuI.pe._201_ AuI.pe._372_ AuI.pe._373_ AuI.pe._101_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._208_ sky130_fd_sc_hd__or4_2
XFILLER_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4729_ MuI._0444_ vssd1 vssd1 vccd1 vccd1 MuI._0445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11331__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _02237_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__nor2_1
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06835_ net58 vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__clkbuf_4
XAuI.pe._589_ AuI.pe._141_ AuI.pe._143_ AuI.pe._074_ vssd1 vssd1 vccd1 vccd1 AuI.pe._144_
+ sky130_fd_sc_hd__a21o_1
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09554_ _02183_ _02184_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__and2b_1
X_06766_ _02905_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__buf_4
XANTENNA__09541__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13084__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07342__A _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__B1 _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _01120_ _01065_ _01122_ _00871_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__a211oi_1
X_06697_ _02118_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__and3_1
X_09485_ _02106_ _02109_ _02108_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a21o_1
XFILLER_211_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08436_ _01007_ _01051_ _01052_ _01053_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a211oi_1
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._140_ FuI._002_ net146 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[11\] sky130_fd_sc_hd__dlxtn_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08367_ _00963_ _00964_ _00969_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__a21o_1
XANTENNA__11398__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__D _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._071_ FuI.a_operand\[28\] FuI.a_operand\[29\] net105 FuI.a_operand\[27\] vssd1
+ vssd1 vccd1 vccd1 FuI._039_ sky130_fd_sc_hd__and4bb_1
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07318_ _06589_ _06592_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__nor2_1
XFILLER_137_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09269__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08173__A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _03335_ _04057_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__nand2_1
XFILLER_109_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08604__C _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._579__B1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__B _04076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _06548_ _05498_ _05563_ _02291_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__a22o_1
XFILLER_192_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _02708_ _02753_ _02945_ _03928_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08901__A _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09763__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10191_ _02861_ _02865_ _02868_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__and4_1
XANTENNA__09716__B _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4259__A2_N MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12901_ _02984_ _05767_ _03257_ _02983_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a22oi_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11873__A2 _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _05636_ _05635_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2b_1
XAuI._1170_ AuI._0367_ AuI._0376_ vssd1 vssd1 vccd1 vccd1 AuI._0377_ sky130_fd_sc_hd__xnor2_1
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09818__A2 _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _05637_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xor2_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08067__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _04510_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _05475_ _05477_ _05564_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._5538__D MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11645_ _04436_ _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__xor2_4
XFILLER_168_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 a_operand[19] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput26 a_operand[29] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_4
X_11576_ _04136_ _04138_ _04298_ _04299_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__a211oi_2
Xinput37 b_operand[0] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
XANTENNA__12317__B _05160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 b_operand[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XANTENNA_MuI._3636__A MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput59 b_operand[2] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10061__B2 AuI.result\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13315_ _06171_ _06172_ _06174_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10527_ _03231_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__nand3_1
XAuI._0954_ net58 net26 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0166_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._5554__C MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0853__B2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ _02741_ _06154_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__nand2_2
X_10458_ _03021_ _03025_ _03022_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21bai_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08811__A _01427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0885_ AuI._0104_ net113 AuI._0098_ vssd1 vssd1 vccd1 vccd1 AuI._0105_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6750_ MuI._2481_ MuI._2667_ vssd1 vssd1 vccd1 vccd1 MuI._2668_ sky130_fd_sc_hd__nor2_1
XMuI._3962_ MuI._3060_ MuI._3061_ vssd1 vssd1 vccd1 vccd1 MuI._3062_ sky130_fd_sc_hd__and2_1
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ FuI.Integer\[24\] _04627_ _02718_ _05595_ _06083_ vssd1 vssd1 vccd1 vccd1
+ _06084_ sky130_fd_sc_hd__a221o_1
XFILLER_112_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10389_ _03081_ _03083_ _03084_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__nand3_1
XMuI._5701_ MuI._1019_ MuI._1022_ vssd1 vssd1 vccd1 vccd1 MuI._1514_ sky130_fd_sc_hd__and2_1
XFILLER_151_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6681_ MuI._0146_ MuI._0787_ MuI._2582_ MuI._0788_ vssd1 vssd1 vccd1 vccd1 MuI._2592_
+ sky130_fd_sc_hd__o31a_1
XFILLER_112_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07427__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3893_ MuI._2988_ MuI._2989_ MuI._2972_ vssd1 vssd1 vccd1 vccd1 MuI._2993_ sky130_fd_sc_hd__a21o_1
X_12128_ _04831_ _04842_ _04844_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__nand3_1
XFILLER_97_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5632_ MuI._1423_ MuI._1437_ vssd1 vssd1 vccd1 vccd1 MuI._1438_ sky130_fd_sc_hd__nor2_1
XAuI._1506_ AuI._0686_ AuI._0687_ AuI._0690_ AuI._0691_ vssd1 vssd1 vccd1 vccd1 AuI._0692_
+ sky130_fd_sc_hd__a31o_2
X_12059_ _02844_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07146__B _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._512_ AuI.pe._071_ vssd1 vssd1 vccd1 vccd1 AuI.pe._072_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5563_ MuI._1313_ MuI._1319_ MuI._1317_ vssd1 vssd1 vccd1 vccd1 MuI._1363_ sky130_fd_sc_hd__a21oi_1
XAuI._1437_ AuI._0503_ AuI._0493_ vssd1 vssd1 vccd1 vccd1 AuI._0623_ sky130_fd_sc_hd__and2_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1030__A1 net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._443_ AuI.pe.significand\[6\] AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1
+ AuI.pe._010_ sky130_fd_sc_hd__nor2_1
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4514_ MuI._0206_ MuI._0208_ vssd1 vssd1 vccd1 vccd1 MuI._0209_ sky130_fd_sc_hd__xor2_1
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5101__B1 MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5494_ MuI._1282_ MuI._1284_ MuI._1233_ MuI._1286_ vssd1 vssd1 vccd1 vccd1 MuI._1287_
+ sky130_fd_sc_hd__a211o_1
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1368_ AuI._0257_ AuI._0558_ AuI._0559_ AuI._0560_ vssd1 vssd1 vccd1 vccd1 AuI._0561_
+ sky130_fd_sc_hd__nand4_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4445_ MuI._3239_ MuI._3359_ MuI._3366_ MuI._3375_ vssd1 vssd1 vccd1 vccd1 MuI._0133_
+ sky130_fd_sc_hd__o31a_1
XANTENNA__07162__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1299_ AuI._0496_ AuI._0497_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[13\]
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4376_ MuI._3326_ MuI._0057_ vssd1 vssd1 vccd1 vccd1 MuI._0058_ sky130_fd_sc_hd__xnor2_1
X_09270_ _01885_ _01886_ _01887_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o21bai_1
XFILLER_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5404__A1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6115_ MuI._1966_ MuI._1969_ vssd1 vssd1 vccd1 vccd1 MuI._1970_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._5404__B2 MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08221_ _00836_ _00838_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3966__A1 MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6046_ MuI._1483_ MuI._2583_ vssd1 vssd1 vccd1 vccd1 MuI._1894_ sky130_fd_sc_hd__nand2_1
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _00768_ _00769_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__and2_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09442__B1 _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _06415_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08083_ _00698_ _00699_ _00700_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__a21o_1
XFILLER_147_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout115_A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ _05788_ _02042_ _02151_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__and3_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11001__B1 _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._448__B AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12243__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6879_ MuI.b_operand\[31\] MuI.a_operand\[31\] vssd1 vssd1 vccd1 vccd1 MuI._2777_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07220__A2 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _01467_ _01461_ _01466_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__nand3_1
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07936_ _00549_ _00552_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3712__C MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11855__A2 _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07867_ _00347_ _00348_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__nand2_1
XFILLER_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _02240_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__xnor2_1
X_06818_ _03465_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[25\] sky130_fd_sc_hd__clkbuf_1
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07798_ _00411_ _00413_ _00415_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__or3_1
XANTENNA__08168__A _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07072__A _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ _02079_ _02167_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__nor2_1
XANTENNA__11306__B _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _02723_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__and3_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _06494_ _00150_ net6 net7 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__and4_1
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _01020_ _01021_ _01019_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__o21bai_1
XFILLER_196_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._123_ FuI._052_ FuI._056_ FuI._024_ FuI.a_operand\[18\] vssd1 vssd1 vccd1 vccd1
+ FuI._008_ sky130_fd_sc_hd__o31a_1
X_09399_ _01996_ _02014_ _02015_ _02016_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__and4_1
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3957__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08615__B _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _04204_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08236__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B2 _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1088__A1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11361_ _04129_ _04130_ _03893_ _04114_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__a211o_1
XANTENNA__11041__B _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10594__A2 _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0835__B2 net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13100_ _04678_ _05929_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__nand2_1
X_10312_ _02958_ _03001_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__xor2_2
XANTENNA_MuI._6189__D MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ _00063_ _00062_ _05445_ _05509_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand4_1
XANTENNA__11976__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ _02715_ _02714_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a21oi_1
X_13031_ _04677_ _05847_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__and2_1
XANTENNA__13249__A _06157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6659__B1 MuI._2559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11543__B2 AuI.result\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10174_ _03067_ _05134_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
XANTENNA_input45_A b_operand[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13296__A1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12099__A2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1012__A1 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10219__A_N _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12299__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6706__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1222_ AuI._0420_ AuI._0425_ vssd1 vssd1 vccd1 vccd1 AuI._0426_ sky130_fd_sc_hd__nor2_1
XFILLER_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1153_ net31 net63 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0361_ sky130_fd_sc_hd__mux2_1
X_12815_ _05608_ _05609_ _05497_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a21boi_1
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07413__C _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4230_ MuI._3200_ MuI._3199_ vssd1 vssd1 vccd1 vccd1 MuI._3330_ sky130_fd_sc_hd__nor2_1
XFILLER_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ _05618_ _05619_ _05615_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a21o_1
XAuI._1084_ AuI._0290_ AuI._0291_ AuI._0293_ AuI._0294_ AuI._0274_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0295_ sky130_fd_sc_hd__mux4_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08806__A _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4161_ MuI._3259_ MuI._3260_ vssd1 vssd1 vccd1 vccd1 MuI._3261_ sky130_fd_sc_hd__nor2_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12677_ _05545_ _05546_ _05527_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4092_ MuI._1472_ MuI._2867_ MuI._2869_ MuI._1010_ vssd1 vssd1 vccd1 vccd1 MuI._3192_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _04385_ _04244_ _04418_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211a_2
XFILLER_30_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _04344_ _02890_ _02928_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07986__B1 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._549__A AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0937_ AuI._0148_ AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 AuI._0149_ sky130_fd_sc_hd__or2b_1
XFILLER_171_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6802_ MuI._2722_ MuI._2723_ MuI._2724_ vssd1 vssd1 vccd1 vccd1 MuI._2725_ sky130_fd_sc_hd__and3_1
XFILLER_171_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4994_ MuI._0725_ MuI._0734_ MuI._0709_ MuI._0736_ vssd1 vssd1 vccd1 vccd1 MuI._0737_
+ sky130_fd_sc_hd__o211ai_4
X_13229_ _06055_ _06101_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__o21a_1
XANTENNA__08898__D _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0868_ AuI._0087_ AuI._0084_ AuI._0079_ vssd1 vssd1 vccd1 vccd1 AuI._0088_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3945_ MuI._2973_ MuI._2977_ MuI._2974_ vssd1 vssd1 vccd1 vccd1 MuI._3045_ sky130_fd_sc_hd__o21bai_1
XMuI._6733_ MuI._2444_ MuI._2648_ vssd1 vssd1 vccd1 vccd1 MuI._2650_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07157__A _06452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6114__A2 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4125__B2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6664_ MuI._0550_ MuI._2573_ vssd1 vssd1 vccd1 vccd1 MuI._2574_ sky130_fd_sc_hd__xor2_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3876_ MuI._2838_ vssd1 vssd1 vccd1 vccd1 MuI._2976_ sky130_fd_sc_hd__clkbuf_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ _01382_ _01387_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__or2b_1
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06996__A _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5615_ MuI._1386_ MuI._1419_ vssd1 vssd1 vccd1 vccd1 MuI._1420_ sky130_fd_sc_hd__xnor2_1
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07313__A1_N _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6595_ MuI._0240_ MuI._2496_ MuI._2497_ vssd1 vssd1 vccd1 vccd1 MuI._2498_ sky130_fd_sc_hd__a21o_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07721_ _00335_ _00336_ _00338_ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__or3_2
XANTENNA__11837__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12510__B _02584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5546_ MuI._1311_ MuI._1302_ MuI._1310_ vssd1 vssd1 vccd1 vccd1 MuI._1344_ sky130_fd_sc_hd__nand3_1
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11407__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13039__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ net114 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__buf_4
XANTENNA__10311__A _02977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._426_ AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 AuI.pe._393_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5477_ MuI._1243_ MuI._1244_ MuI._1259_ vssd1 vssd1 vccd1 vccd1 MuI._1268_ sky130_fd_sc_hd__a21o_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _00198_ _00200_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__xor2_1
XFILLER_81_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11126__B _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__C _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4428_ MuI._0109_ MuI._0113_ vssd1 vssd1 vccd1 vccd1 MuI._0114_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12798__B1 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _01895_ _01889_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__or2b_1
XFILLER_40_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1367__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4359_ MuI._2840_ MuI._2867_ MuI._2869_ MuI._2843_ vssd1 vssd1 vccd1 vccd1 MuI._0039_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._5756__A MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _01203_ _01211_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__nand2_1
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _00820_ _00821_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__nor2_1
X_09184_ _00877_ _00011_ _06446_ _04111_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._5475__B MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12014__A2 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6029_ MuI._1873_ MuI._1874_ vssd1 vssd1 vccd1 vccd1 MuI._1875_ sky130_fd_sc_hd__nor2_1
X_08135_ _00751_ _00752_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__nor2_1
XFILLER_175_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07977__B1 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _00682_ _00683_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07017_ _05606_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[25\] sky130_fd_sc_hd__buf_4
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10205__B _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08968_ _01528_ _01530_ _01584_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a211o_1
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4667__A2 MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07919_ _06564_ _02474_ _05101_ _05176_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__and4_1
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4835__A MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ _06593_ _04520_ _01514_ _01515_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12420__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ _03660_ _03665_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__or2_1
XFILLER_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09432__D _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _03589_ _03590_ _03437_ _03439_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__o211a_1
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _05462_ _05463_ _05289_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__o21ai_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _03733_ _04251_ _03348_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__nand3_1
XFILLER_158_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10875__B _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _03024_ _02721_ _02853_ _04011_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__a22o_1
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6041__A1 MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _05314_ _05315_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13202__A1 _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._106_ FuI._037_ net104 FuI._056_ vssd1 vssd1 vccd1 vccd1 FuI._063_ sky130_fd_sc_hd__and3b_1
XANTENNA__13202__B2 _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ _04029_ _04032_ _04030_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__o21bai_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0808__A1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ _05242_ _05136_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__nor2_1
XFILLER_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11344_ _03721_ _03726_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07432__A2 _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__A1 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1306__A AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11275_ _04034_ _04036_ _04037_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12713__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__A2 _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ _05822_ _05865_ _05907_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__or3_1
X_10226_ _02781_ _02909_ _02780_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a21o_1
XMuI._3730_ MuI._2829_ vssd1 vssd1 vccd1 vccd1 MuI._2830_ sky130_fd_sc_hd__clkbuf_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10157_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__inv_2
XFILLER_94_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3661_ MuI._2616_ vssd1 vssd1 vccd1 vccd1 MuI._2627_ sky130_fd_sc_hd__buf_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _02345_ _04186_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__and2b_1
XMuI._5400_ MuI._1119_ MuI._1171_ vssd1 vssd1 vccd1 vccd1 MuI._1183_ sky130_fd_sc_hd__xnor2_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6380_ MuI._2789_ MuI._0438_ vssd1 vssd1 vccd1 vccd1 MuI._2261_ sky130_fd_sc_hd__nand2_1
XMuI._3592_ MuI._0350_ MuI._1285_ MuI._1318_ MuI._0526_ vssd1 vssd1 vccd1 vccd1 MuI._1868_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10131__A _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5331_ MuI._1101_ MuI._1104_ MuI._1105_ MuI._1106_ vssd1 vssd1 vccd1 vccd1 MuI._1107_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1205_ AuI._0262_ AuI._0330_ AuI._0274_ AuI._0294_ vssd1 vssd1 vccd1 vccd1 AuI._0410_
+ sky130_fd_sc_hd__or4b_1
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5262_ MuI._0327_ MuI._0477_ MuI._3306_ MuI._3307_ vssd1 vssd1 vccd1 vccd1 MuI._1031_
+ sky130_fd_sc_hd__and4_1
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._551__B AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1136_ AuI._0344_ vssd1 vssd1 vccd1 vccd1 AuI._0345_ sky130_fd_sc_hd__inv_2
XFILLER_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4213_ MuI._2843_ MuI._2871_ vssd1 vssd1 vccd1 vccd1 MuI._3313_ sky130_fd_sc_hd__nand2_1
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07440__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5193_ MuI._0855_ MuI._0854_ MuI._0853_ vssd1 vssd1 vccd1 vccd1 MuI._0956_ sky130_fd_sc_hd__o21ai_1
XFILLER_204_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _00125_ _05884_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__nand2_1
XAuI._1067_ net64 net124 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0278_ sky130_fd_sc_hd__mux2_1
XANTENNA_MuI._4480__A MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__D _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4144_ MuI._3242_ MuI._3243_ vssd1 vssd1 vccd1 vccd1 MuI._3244_ sky130_fd_sc_hd__nor2_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4075_ MuI._3172_ MuI._3173_ MuI._3174_ vssd1 vssd1 vccd1 vccd1 MuI._3175_ sky130_fd_sc_hd__a21oi_1
XFILLER_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5543__B1 MuI._2876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09940_ _02588_ _02589_ _02328_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09086__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4977_ MuI._1296_ MuI._1791_ MuI.a_operand\[3\] MuI._0444_ vssd1 vssd1 vccd1
+ vccd1 MuI._0718_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3543__B MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09871_ _02501_ _02508_ _02510_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a21oi_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1224__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12180__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6716_ MuI._2621_ MuI._2626_ MuI._2630_ vssd1 vssd1 vccd1 vccd1 MuI._2631_ sky130_fd_sc_hd__and3_1
XMuI._3928_ MuI._2995_ MuI._3026_ vssd1 vssd1 vccd1 vccd1 MuI._3028_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08822_ _00150_ net14 _05176_ _06494_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a22oi_2
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__A2 _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6647_ MuI._2554_ MuI._2523_ vssd1 vssd1 vccd1 vccd1 MuI._2555_ sky130_fd_sc_hd__xnor2_1
XMuI._3859_ MuI._2956_ MuI._2949_ MuI._2955_ vssd1 vssd1 vccd1 vccd1 MuI._2959_ sky130_fd_sc_hd__o21ai_1
X_08753_ _01356_ _01370_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__nor2_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07704_ net113 net54 _04165_ _00266_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__and4_1
XMuI._6578_ MuI._0548_ MuI._2478_ MuI._0988_ MuI._0691_ vssd1 vssd1 vccd1 vccd1 MuI._2479_
+ sky130_fd_sc_hd__and4b_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08684_ _01017_ _01018_ _01048_ _01049_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5529_ MuI._1316_ MuI._1314_ vssd1 vssd1 vccd1 vccd1 MuI._1325_ sky130_fd_sc_hd__and2b_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07635_ _00212_ _00213_ _00251_ _00252_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__a22oi_2
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__B1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5074__A2 MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._409_ AuI.pe.significand\[3\] AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1
+ AuI.pe._376_ sky130_fd_sc_hd__or2b_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._467__A2 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07566_ _00171_ _00172_ _00183_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13432__B2 _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09305_ _01921_ _01922_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nor2_1
XANTENNA__10246__A1 _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07350__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07497_ _00112_ _00113_ _00114_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__nand3_1
XFILLER_139_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09236_ _01298_ _01299_ _01242_ _01300_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__or4bb_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4585__A1 MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4585__B2 MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09167_ _01714_ _01716_ _01715_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__o21ai_1
XFILLER_163_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _00088_ _00040_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__nand2_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _02647_ _00592_ _00089_ _02582_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a22oi_2
XANTENNA__11957__D _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08049_ _00483_ _00519_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__or2_1
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4549__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__D net123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__xnor2_1
XFILLER_150_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _02677_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__and2_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10721__A2 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0974__A0 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__C net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11962_ _04775_ _04776_ _04771_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a21o_1
XFILLER_44_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _03377_ _03474_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__a21oi_2
XFILLER_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4715__D MuI._0228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11893_ _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nand2_1
XFILLER_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10844_ _00124_ _00125_ _06603_ _06605_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__and4_1
XFILLER_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07260__A _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10775_ _03489_ _03491_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__a21o_1
XFILLER_201_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4731__C MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12514_ _02800_ _05255_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o21ai_1
XFILLER_185_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13494_ _06408_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_145_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _05296_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__xnor2_1
XFILLER_166_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__A _00707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _05222_ _05223_ _05181_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__o21a_1
XMuI._4900_ MuI._0632_ vssd1 vssd1 vccd1 vccd1 MuI._0633_ sky130_fd_sc_hd__inv_2
XMuI._5880_ MuI._1647_ MuI._1710_ vssd1 vssd1 vccd1 vccd1 MuI._1711_ sky130_fd_sc_hd__xnor2_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11327_ _04092_ _04093_ _04026_ _04027_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o211ai_4
XANTENNA_MuI._6020__A MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10126__A _02801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4831_ MuI._2843_ MuI._3268_ MuI._0503_ MuI._0505_ vssd1 vssd1 vccd1 vccd1 MuI._0557_
+ sky130_fd_sc_hd__o2bb2a_1
XAuI.pe._760_ AuI.pe._071_ AuI.pe._197_ AuI.pe._397_ vssd1 vssd1 vccd1 vccd1 AuI.pe._304_
+ sky130_fd_sc_hd__a21o_1
XANTENNA__10960__A2 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output76_A net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _02750_ _03855_ _03856_ _04010_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__a311o_1
XFILLER_68_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12162__A1 _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4762_ MuI._0478_ MuI._0480_ vssd1 vssd1 vccd1 vccd1 MuI._0481_ sky130_fd_sc_hd__nor2_1
XAuI.pe._691_ AuI.pe._211_ AuI.pe._208_ AuI.pe._385_ vssd1 vssd1 vccd1 vccd1 AuI.pe._239_
+ sky130_fd_sc_hd__o21ai_1
X_10209_ _02787_ _02890_ _02789_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08905__A2 _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ _03771_ _03754_ _03756_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__nand3_2
XMuI._3713_ MuI._2811_ vssd1 vssd1 vccd1 vccd1 MuI._2813_ sky130_fd_sc_hd__buf_2
XMuI._6501_ MuI._2393_ MuI._2001_ MuI._1995_ vssd1 vssd1 vccd1 vccd1 MuI._2394_ sky130_fd_sc_hd__a21oi_1
XFILLER_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4693_ MuI._0401_ MuI._0402_ vssd1 vssd1 vccd1 vccd1 MuI._0406_ sky130_fd_sc_hd__nor2_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6432_ MuI._2315_ MuI._2316_ MuI._2317_ vssd1 vssd1 vccd1 vccd1 MuI._2318_ sky130_fd_sc_hd__or3_1
XMuI._3644_ MuI._2429_ vssd1 vssd1 vccd1 vccd1 MuI._2440_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10499__C _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4906__C MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09072__D net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12995__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6363_ MuI._2197_ MuI._2195_ vssd1 vssd1 vccd1 vccd1 MuI._2243_ sky130_fd_sc_hd__xor2_1
XANTENNA_AuI.pe._562__A AuI.pe.significand\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3575_ MuI._1131_ MuI._1219_ MuI._1560_ MuI._1670_ vssd1 vssd1 vccd1 vccd1 MuI._1681_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._4625__D MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5314_ MuI._2895_ MuI._0101_ vssd1 vssd1 vccd1 vccd1 MuI._1089_ sky130_fd_sc_hd__nand2_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6253__B2 MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__A _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6294_ MuI._2163_ MuI._2166_ vssd1 vssd1 vccd1 vccd1 MuI._2167_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07420_ net40 net41 _06611_ _06602_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__and4_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4264__B1 MuI._3363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08266__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5245_ MuI._0939_ MuI._0945_ MuI._1012_ vssd1 vssd1 vccd1 vccd1 MuI._1013_ sky130_fd_sc_hd__a21o_1
XFILLER_204_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1119_ AuI._0322_ AuI._0323_ vssd1 vssd1 vccd1 vccd1 AuI._0328_ sky130_fd_sc_hd__and2_1
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3819__A MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ _06479_ _06480_ _06461_ _05627_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__and4_1
XANTENNA__07601__C _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5176_ MuI._0932_ MuI._0936_ vssd1 vssd1 vccd1 vccd1 MuI._0937_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ net38 vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__buf_4
XMuI._4127_ MuI._1285_ MuI._2363_ MuI._3226_ MuI._3224_ vssd1 vssd1 vccd1 vccd1 MuI._3227_
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13178__B1 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ _01635_ _01636_ _01637_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4360__D MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13111__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4058_ MuI._3082_ MuI._3083_ vssd1 vssd1 vccd1 vccd1 MuI._3158_ sky130_fd_sc_hd__xor2_2
XANTENNA__11728__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09097__A net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10036__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09923_ _02402_ _02447_ _02583_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__and3b_2
XFILLER_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3704__D MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09854_ _02458_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07990__D _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08805_ _01419_ _01422_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__or2b_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__B2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13066__B _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ _02366_ _02373_ _02372_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__o21a_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5295__A2 MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06997_ _05391_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__clkbuf_4
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _02582_ _02647_ _00082_ _00084_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3720__C MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09560__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _01279_ _01280_ _01284_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a21o_1
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07618_ _03152_ _00047_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__and2_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _02485_ _04832_ _04896_ _06565_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a22oi_1
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07080__A _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09085__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _00160_ _00166_ vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09085__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _03080_ _03267_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08832__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08832__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _01832_ _01835_ _01836_ _01732_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a211oi_2
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10491_ _03192_ _03193_ _03194_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nand3_1
XANTENNA__12426__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12916__B1 _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__A _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__inv_2
XFILLER_182_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08342__C net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3464__A MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _04902_ _04903_ _04991_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a211oi_2
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _03731_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__inv_2
XANTENNA__08061__D _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12092_ _00727_ _06546_ _03051_ _00728_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22oi_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08348__B1 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4730__A1 MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4730__B2 MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1470_ AuI._0320_ AuI._0323_ vssd1 vssd1 vccd1 vccd1 AuI._0656_ sky130_fd_sc_hd__and2_1
X_11043_ _03786_ _03787_ _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__or3_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _05885_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _04759_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nand2b_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6786__A2 MuI._2563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11876_ _04684_ _04685_ _04686_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__or3_1
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3639__A MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10827_ _03534_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5030_ MuI._0771_ MuI._0775_ vssd1 vssd1 vccd1 vccd1 MuI._0776_ sky130_fd_sc_hd__and2_2
XANTENNA_MuI._4461__C MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__A1 _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11958__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1675__A1 net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _03137_ _03480_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a21oi_4
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__A2_N _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13477_ _01328_ _01329_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nor2_1
X_10689_ _03404_ _03405_ _03406_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a21o_1
XANTENNA__08533__B _01150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _05276_ _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__o21ai_1
XFILLER_127_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5932_ MuI._1716_ MuI._1755_ MuI._1767_ vssd1 vssd1 vccd1 vccd1 MuI._1768_ sky130_fd_sc_hd__a21bo_1
XFILLER_126_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12359_ _06439_ _05123_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nand2_1
XANTENNA__07149__B _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._812_ AuI.pe.significand\[10\] AuI.pe.significand\[11\] AuI.pe.significand\[12\]
+ AuI.pe.significand\[9\] vssd1 vssd1 vccd1 vccd1 AuI.pe._351_ sky130_fd_sc_hd__or4b_1
XFILLER_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5863_ MuI._0685_ MuI._1691_ vssd1 vssd1 vccd1 vccd1 MuI._1693_ sky130_fd_sc_hd__nor2_1
XFILLER_141_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11894__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._743_ AuI.pe._120_ AuI.pe._079_ AuI.pe._285_ AuI.pe._386_ AuI.pe._287_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._288_ sky130_fd_sc_hd__a221o_1
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4814_ MuI._0536_ MuI._0538_ vssd1 vssd1 vccd1 vccd1 MuI._0539_ sky130_fd_sc_hd__xnor2_1
X_06920_ net6 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__clkbuf_4
XMuI._5794_ MuI._2660_ MuI._2429_ MuI._3306_ MuI._2880_ vssd1 vssd1 vccd1 vccd1 MuI._1617_
+ sky130_fd_sc_hd__and4_1
XAuI._1668_ AuI.exponent_sub\[6\] AuI._0599_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0020_
+ sky130_fd_sc_hd__o21a_1
XFILLER_110_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._674_ AuI.pe._102_ AuI.pe._112_ AuI.pe._079_ AuI.pe._142_ AuI.pe._222_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._223_ sky130_fd_sc_hd__a221o_1
XANTENNA__07165__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4745_ MuI._0353_ MuI._0352_ vssd1 vssd1 vccd1 vccd1 MuI._0463_ sky130_fd_sc_hd__nor2_1
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06851_ _03820_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1599_ AuI._0626_ AuI._0766_ AuI._0621_ vssd1 vssd1 vccd1 vccd1 AuI._0771_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4676_ MuI._0343_ MuI._0345_ vssd1 vssd1 vccd1 vccd1 MuI._0387_ sky130_fd_sc_hd__and2_1
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09570_ _02193_ _02201_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a21bo_1
X_06782_ _03078_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6415_ MuI._2296_ MuI._2299_ vssd1 vssd1 vccd1 vccd1 MuI._2300_ sky130_fd_sc_hd__and2b_1
XMuI._3627_ MuI._1560_ MuI._2242_ vssd1 vssd1 vccd1 vccd1 MuI._2253_ sky130_fd_sc_hd__nor2_1
XFILLER_209_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ _01096_ _01103_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__and2_1
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08708__B _01325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3558_ MuI._1483_ vssd1 vssd1 vccd1 vccd1 MuI._1494_ sky130_fd_sc_hd__clkbuf_4
XMuI._6346_ MuI._2217_ MuI._2223_ vssd1 vssd1 vccd1 vccd1 MuI._2224_ sky130_fd_sc_hd__nand2_1
XANTENNA__11415__A _02905_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07612__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _00886_ _01068_ _01069_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._5748__B MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6277_ MuI._2056_ MuI._2061_ MuI._2147_ vssd1 vssd1 vccd1 vccd1 MuI._2148_ sky130_fd_sc_hd__a21oi_1
X_07403_ _06678_ _06679_ _00019_ _00020_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__o211ai_2
XFILLER_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._3489_ MuI.b_operand\[19\] vssd1 vssd1 vccd1 vccd1 MuI._0735_ sky130_fd_sc_hd__buf_2
XANTENNA_MuI._3549__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__B _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08383_ _00999_ _01000_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__and2b_1
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5228_ MuI._0904_ MuI._0903_ vssd1 vssd1 vccd1 vccd1 MuI._0994_ sky130_fd_sc_hd__or2b_1
XANTENNA__11949__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12071__B1 _04891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ _06629_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__xnor2_2
XFILLER_177_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5159_ MuI._0915_ MuI._0916_ MuI._0914_ vssd1 vssd1 vccd1 vccd1 MuI._0918_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5764__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _06565_ _02485_ _06562_ _06476_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__nand4_1
XFILLER_136_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09004_ _01590_ _01591_ _01618_ _01621_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__o211ai_1
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ _06490_ _06493_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o21bai_1
XFILLER_118_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11392__A1_N _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09906_ _02545_ _02553_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__nand3_1
XFILLER_120_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09274__B _01891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__A_N _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0929__B1 net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3731__B MuI._0449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _02438_ _02480_ _02477_ _02479_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09542__A2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11309__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5848__A2_N MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ net111 net126 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__nand2_1
XFILLER_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09290__A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4265__D MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08719_ _02528_ _04585_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__nand2_1
XANTENNA__07803__A _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _02319_ _02321_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__or2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11970__D _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1354__B1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _03324_ _05198_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__nand2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _04452_ _04453_ _04449_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a21o_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _04161_ _06302_ _06303_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__a31o_1
XFILLER_211_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ _02767_ _02882_ _02884_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__a21o_1
XFILLER_211_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11592_ _04230_ _04366_ _04379_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o21a_1
XFILLER_195_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5096__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5674__A MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13331_ _06239_ _06240_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__and2_1
XFILLER_167_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10543_ _03245_ _03249_ _03251_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__nand3_1
XFILLER_195_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0970_ AuI._0164_ AuI._0169_ AuI._0181_ vssd1 vssd1 vccd1 vccd1 AuI._0182_ sky130_fd_sc_hd__and3_1
XANTENNA__09094__A2_N _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13262_ _06168_ _06169_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a21boi_1
XANTENNA_AuI.pe._597__B2 AuI.pe._089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _03175_ _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12213_ _04769_ _04912_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2b_1
XFILLER_136_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _02837_ _06097_ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__o21a_1
XFILLER_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__B1 _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09465__A _02069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _04957_ _04847_ _04973_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a211o_1
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08800__C _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1522_ AuI.pe.Significand\[1\] AuI._0695_ vssd1 vssd1 vccd1 vccd1 AuI._0707_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__B _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _04899_ _02896_ _02928_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__mux2_1
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ _03761_ _03770_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__xor2_2
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1453_ AuI._0451_ AuI._0454_ vssd1 vssd1 vccd1 vccd1 AuI._0639_ sky130_fd_sc_hd__xnor2_2
XMuI._4530_ MuI._0215_ MuI._0223_ MuI._0225_ vssd1 vssd1 vccd1 vccd1 MuI._0226_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10123__B _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4467__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1384_ AuI._0375_ AuI._0498_ AuI._0574_ vssd1 vssd1 vccd1 vccd1 AuI._0575_ sky130_fd_sc_hd__or3_1
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4461_ MuI.a_operand\[21\] MuI.a_operand\[20\] MuI.b_operand\[1\] MuI.b_operand\[0\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0150_ sky130_fd_sc_hd__and4_1
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._521__A1 AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._521__B2 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12977_ _02980_ _03444_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__and2_1
XFILLER_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6200_ MuI._2043_ MuI._2045_ MuI._2062_ vssd1 vssd1 vccd1 vccd1 MuI._2063_ sky130_fd_sc_hd__or3_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4392_ MuI._0051_ MuI._0073_ MuI._0074_ vssd1 vssd1 vccd1 vccd1 MuI._0075_ sky130_fd_sc_hd__a21oi_2
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11928_ _04740_ _04741_ _04721_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__a21o_1
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6131_ MuI._1849_ MuI._1907_ vssd1 vssd1 vccd1 vccd1 MuI._1987_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._4472__B MuI._0154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ _04663_ _04666_ _04667_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__nand3_1
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13481__A1_N _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6062_ MuI._3033_ MuI._1910_ vssd1 vssd1 vccd1 vccd1 MuI._1911_ sky130_fd_sc_hd__nor2_1
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5013_ MuI._0755_ MuI._0756_ vssd1 vssd1 vccd1 vccd1 MuI._0758_ sky130_fd_sc_hd__and2b_1
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3519__D MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5584__A MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07050_ _05959_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._5195__B2 MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12356__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0871__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12356__B2 _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 Underflow sky130_fd_sc_hd__buf_2
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5915_ MuI._1746_ MuI._1748_ MuI._1741_ MuI._1742_ vssd1 vssd1 vccd1 vccd1 MuI._1750_
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12513__B _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12108__A1 _04803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5846_ MuI._1576_ MuI._1578_ vssd1 vssd1 vccd1 vccd1 MuI._1674_ sky130_fd_sc_hd__nand2_1
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07952_ _00567_ _00569_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__nand2_1
XFILLER_130_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._726_ AuI.pe._270_ AuI.pe._271_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._272_
+ sky130_fd_sc_hd__a21o_1
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06903_ _04380_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__clkbuf_4
XMuI._5777_ MuI._1520_ MuI._1523_ MuI._1521_ vssd1 vssd1 vccd1 vccd1 MuI._1598_ sky130_fd_sc_hd__o21ba_1
X_07883_ _00499_ _00500_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__xnor2_2
XFILLER_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._657_ AuI.pe._046_ AuI.pe._164_ AuI.pe._397_ AuI.pe._028_ AuI.pe._206_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._207_ sky130_fd_sc_hd__a221o_1
XANTENNA__11331__A2 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4728_ MuI.a_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._0444_ sky130_fd_sc_hd__buf_2
X_09622_ _02226_ _02234_ _02236_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__and3_1
X_06834_ _03637_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[28\] sky130_fd_sc_hd__clkbuf_1
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08719__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._588_ AuI.pe._106_ AuI.pe._125_ AuI.pe._101_ AuI.pe._142_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._143_ sky130_fd_sc_hd__o31ai_1
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4659_ MuI._0366_ MuI._0364_ vssd1 vssd1 vccd1 vccd1 MuI._0368_ sky130_fd_sc_hd__and2b_1
X_09553_ _02183_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09541__C _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06765_ _02894_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13084__A2 _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ _00868_ _00869_ _01121_ _00849_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07342__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__B2 AuI.result\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _02106_ _02108_ _02109_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__nand3_1
X_06696_ _02151_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._750__A AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6329_ MuI._2185_ MuI._2204_ vssd1 vssd1 vccd1 vccd1 MuI._2205_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08435_ _00835_ _00844_ _00845_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__and3_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ _00977_ _00982_ _00983_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08454__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFuI._070_ net104 vssd1 vssd1 vccd1 vccd1 FuI._038_ sky130_fd_sc_hd__inv_2
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08799__B1 _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ _06523_ _06531_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__or2b_1
XANTENNA__09269__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08297_ _00911_ _00914_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__and2b_2
XANTENNA__08173__B net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._579__A1 AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _02291_ _06548_ _05498_ _06461_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__and4_1
XANTENNA__08604__D _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10358__B1 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ net109 vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__buf_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08901__B _01350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09285__A _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nor2_2
XFILLER_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06702__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09716__C _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3742__A MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12900_ _05712_ _05730_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__and2_1
XFILLER_101_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07533__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12831_ _05710_ _05711_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__xnor2_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12762_ _06429_ _05327_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nand2_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ _04371_ _04500_ _04508_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__and3_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10833__A1 _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05475_ _05477_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11644_ _03525_ _04660_ _04256_ _04255_ _04800_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a32o_2
XFILLER_202_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 a_operand[1] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
X_11575_ _03831_ _04542_ _04267_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__nand3_1
Xinput27 a_operand[2] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_4
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 b_operand[10] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_6
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13314_ _06128_ _06191_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__nand2_1
Xinput49 b_operand[20] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_6
XFILLER_183_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _03054_ _03052_ _03053_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a21bo_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0953_ AuI._0110_ AuI._0157_ AuI._0159_ AuI._0161_ AuI._0154_ vssd1 vssd1 vccd1
+ vccd1 AuI._0165_ sky130_fd_sc_hd__a311o_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0853__A2 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__B _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13245_ _02692_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10457_ _03026_ _03034_ _03033_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__a21o_1
XAuI._0884_ net21 vssd1 vssd1 vccd1 vccd1 AuI._0104_ sky130_fd_sc_hd__inv_2
XMuI._3961_ MuI._3053_ MuI._3054_ MuI._3038_ MuI._3059_ vssd1 vssd1 vccd1 vccd1 MuI._3061_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _05531_ _02726_ _02730_ AuI.result\[24\] vssd1 vssd1 vccd1 vccd1 _06083_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13429__B _06305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ _03081_ _03083_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a21o_1
XMuI._5700_ MuI._1510_ MuI._1511_ MuI._1506_ vssd1 vssd1 vccd1 vccd1 MuI._1513_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3892_ MuI._2972_ MuI._2988_ MuI._2989_ vssd1 vssd1 vccd1 vccd1 MuI._2992_ sky130_fd_sc_hd__nand3_1
XMuI._6680_ MuI._2585_ MuI._2590_ MuI._2485_ vssd1 vssd1 vccd1 vccd1 MuI._2591_ sky130_fd_sc_hd__mux2_1
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12127_ _04954_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07427__B _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5631_ MuI._1421_ MuI._1422_ MuI._1380_ vssd1 vssd1 vccd1 vccd1 MuI._1437_ sky130_fd_sc_hd__o21a_1
XAuI._1505_ AuI._0596_ AuI._0688_ AuI._0598_ vssd1 vssd1 vccd1 vccd1 AuI._0691_ sky130_fd_sc_hd__a21bo_1
XFILLER_96_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12058_ _02871_ _04647_ _01233_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o21a_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._511_ AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 AuI.pe._071_ sky130_fd_sc_hd__buf_2
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07146__C _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5562_ MuI._1313_ MuI._1317_ MuI._1319_ vssd1 vssd1 vccd1 vccd1 MuI._1361_ sky130_fd_sc_hd__and3_1
X_11009_ _03750_ _03748_ _03749_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nand3_2
XAuI._1436_ AuI._0515_ AuI._0519_ AuI._0621_ vssd1 vssd1 vccd1 vccd1 AuI._0622_ sky130_fd_sc_hd__o21a_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1030__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._442_ AuI.pe._372_ AuI.pe._394_ AuI.pe._008_ vssd1 vssd1 vccd1 vccd1 AuI.pe._009_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__10521__B1 _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4513_ MuI._0051_ MuI._0073_ vssd1 vssd1 vccd1 vccd1 MuI._0208_ sky130_fd_sc_hd__xor2_2
XFILLER_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5493_ MuI._1231_ MuI._1232_ MuI._1223_ vssd1 vssd1 vccd1 vccd1 MuI._1286_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07443__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1367_ net15 net47 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0560_ sky130_fd_sc_hd__mux2_2
XFILLER_92_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4444_ MuI._0120_ MuI._0124_ MuI._0123_ vssd1 vssd1 vccd1 vccd1 MuI._0132_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1298_ AuI._0484_ AuI._0485_ AuI._0494_ AuI._0495_ vssd1 vssd1 vccd1 vccd1 AuI._0497_
+ sky130_fd_sc_hd__or4_1
XMuI._4375_ MuI._3328_ MuI._3327_ vssd1 vssd1 vccd1 vccd1 MuI._0057_ sky130_fd_sc_hd__nor2_1
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5404__A2 MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6114_ MuI._0581_ MuI._2851_ MuI._1889_ MuI._1968_ vssd1 vssd1 vccd1 vccd1 MuI._1969_
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _00539_ _00837_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__nor2_1
XFILLER_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6045_ MuI._1891_ MuI._1892_ vssd1 vssd1 vccd1 vccd1 MuI._1893_ sky130_fd_sc_hd__xor2_1
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3966__A2 MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _00766_ _00767_ _00419_ _00428_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09442__A1 _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__B1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09442__B2 _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07102_ _05273_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__and2_1
XANTENNA__10166__B_N _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08082_ _00488_ _00490_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__nand2_1
XFILLER_174_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07033_ _05777_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout108_A net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__A1 _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11001__B2 _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._448__C AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12243__B _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6878_ MuI._2504_ MuI._2735_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[30\]
+ sky130_fd_sc_hd__a21oi_1
X_08984_ _01598_ _01600_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a21bo_1
XMuI._5829_ MuI._1263_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._1655_ sky130_fd_sc_hd__nand2_1
X_07935_ _00549_ _00552_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__and2b_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3712__D MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._709_ AuI.pe._393_ AuI.pe._375_ vssd1 vssd1 vccd1 vccd1 AuI.pe._255_ sky130_fd_sc_hd__nor2_1
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07866_ _00235_ _00244_ _00243_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a21o_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ _02377_ _00272_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__nand2_1
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06817_ _03454_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__and3_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07797_ _00414_ _06622_ _05305_ _05370_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__and4_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08168__B _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09536_ _06620_ _03873_ _02077_ _02078_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__o2bb2a_1
X_06748_ _02712_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__buf_6
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13462__C1 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09467_ _02248_ _00098_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__nand2_1
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _00852_ _00854_ _00853_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__o21ai_1
XFILLER_200_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4603__B1 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._122_ FuI._052_ FuI._056_ FuI._024_ FuI._031_ vssd1 vssd1 vccd1 vccd1 FuI._007_
+ sky130_fd_sc_hd__o31a_1
X_09398_ _01994_ _01993_ _01992_ _01981_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__o211ai_1
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3957__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08349_ _06503_ _06504_ _05176_ _05241_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__and4_1
XANTENNA__08236__A2 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _03893_ _04114_ _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__o211ai_2
XANTENNA__11041__C net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0835__A2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10311_ _02977_ _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__xnor2_2
XFILLER_153_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11291_ _00046_ _06666_ _00398_ _00049_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a22o_1
XANTENNA__11976__C _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _01847_ _02639_ _05843_ _03314_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o31a_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10242_ _02926_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__clkbuf_4
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09446__C net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3472__A MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10173_ _02849_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nand2_1
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input38_A b_operand[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10889__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0907__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08172__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__B2 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07263__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1221_ AuI._0422_ AuI._0424_ vssd1 vssd1 vccd1 vccd1 AuI._0425_ sky130_fd_sc_hd__nand2_1
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1152_ AuI._0344_ AuI._0358_ vssd1 vssd1 vccd1 vccd1 AuI._0360_ sky130_fd_sc_hd__nand2_1
XFILLER_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12814_ _05692_ _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__nor2_1
XANTENNA__12256__B1 _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07413__D _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _05615_ _05618_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__nand3_1
XAuI._1083_ AuI._0176_ AuI._0192_ AuI._0198_ vssd1 vssd1 vccd1 vccd1 AuI._0294_ sky130_fd_sc_hd__and3_1
XFILLER_188_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4160_ MuI._3195_ MuI._3188_ MuI._3194_ vssd1 vssd1 vccd1 vccd1 MuI._3260_ sky130_fd_sc_hd__a21oi_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08806__B _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__A _00672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _05527_ _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and3_1
XFILLER_203_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4091_ MuI.a_operand\[19\] MuI._1461_ MuI._3189_ MuI._3190_ vssd1 vssd1 vccd1
+ vccd1 MuI._3191_ sky130_fd_sc_hd__and4_1
XFILLER_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ _04417_ _04398_ _04399_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__nand3_2
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._660__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11558_ _02784_ _04343_ _02785_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__o21bai_1
XANTENNA_AuI._0878__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A1 _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10509_ _03212_ _03195_ _03197_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nand3_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B2 _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0936_ net54 net22 AuI._0121_ vssd1 vssd1 vccd1 vccd1 AuI._0148_ sky130_fd_sc_hd__mux2_1
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _03888_ _03892_ _04127_ _04128_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12344__A _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6801_ MuI._2608_ MuI._2721_ MuI._2687_ vssd1 vssd1 vccd1 vccd1 MuI._2724_ sky130_fd_sc_hd__a21bo_1
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _06134_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and2_1
XMuI._4993_ MuI._0646_ MuI._0708_ MuI._0707_ MuI._0693_ vssd1 vssd1 vccd1 vccd1 MuI._0736_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0867_ AuI._0078_ net6 AuI._0082_ net36 vssd1 vssd1 vccd1 vccd1 AuI._0087_ sky130_fd_sc_hd__o22a_1
XANTENNA_MuI._4478__A MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6732_ MuI._2637_ MuI._2459_ MuI._2469_ vssd1 vssd1 vccd1 vccd1 MuI._2648_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3944_ MuI._3041_ MuI._3042_ MuI._3040_ vssd1 vssd1 vccd1 vccd1 MuI._3044_ sky130_fd_sc_hd__o21ai_1
XFILLER_152_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _05918_ _05988_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__or2_1
XFILLER_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4125__A2 MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6663_ MuI._1837_ MuI._2507_ MuI._0784_ vssd1 vssd1 vccd1 vccd1 MuI._2573_ sky130_fd_sc_hd__a21o_1
XFILLER_112_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3875_ MuI._2853_ vssd1 vssd1 vccd1 vccd1 MuI._2975_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5614_ MuI._1388_ MuI._1387_ vssd1 vssd1 vccd1 vccd1 MuI._1419_ sky130_fd_sc_hd__nor2_1
X_07720_ _06457_ _00337_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__or2_1
XMuI._6594_ MuI._0229_ MuI._0218_ MuI._0196_ vssd1 vssd1 vccd1 vccd1 MuI._2497_ sky130_fd_sc_hd__and3b_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5545_ MuI._1341_ MuI._1342_ vssd1 vssd1 vccd1 vccd1 MuI._1343_ sky130_fd_sc_hd__or2_1
XFILLER_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1419_ AuI._0605_ vssd1 vssd1 vccd1 vccd1 AuI.Exception sky130_fd_sc_hd__dlymetal6s2s_1
X_07651_ _00125_ _00267_ _04305_ _00124_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__a22oi_1
XANTENNA__11407__B _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._425_ AuI.pe.significand\[12\] AuI.pe._388_ AuI.pe._389_ AuI.pe._391_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._392_ sky130_fd_sc_hd__a31o_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._479__B1 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5102__A MuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5476_ MuI._1265_ MuI._1266_ vssd1 vssd1 vccd1 vccd1 MuI._1267_ sky130_fd_sc_hd__xor2_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07582_ _05123_ _00010_ _00199_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__a21bo_1
XANTENNA__07323__D _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4427_ MuI._0112_ MuI._0438_ vssd1 vssd1 vccd1 vccd1 MuI._0113_ sky130_fd_sc_hd__nand2_1
X_09321_ _01926_ _01937_ _01938_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nand3_2
XFILLER_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4358_ MuI._2616_ MuI._2871_ vssd1 vssd1 vccd1 vccd1 MuI._0038_ sky130_fd_sc_hd__nand2_1
X_09252_ _01203_ _01211_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__or2_1
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5756__B MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6586__B1 MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__B1_N _06470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4888__A2_N MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08203_ _06501_ _06548_ _05241_ _06562_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__and4_1
XMuI._4289_ MuI._3340_ MuI._3341_ vssd1 vssd1 vccd1 vccd1 MuI._3389_ sky130_fd_sc_hd__or2b_1
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09183_ _01744_ _01800_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._5475__C MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6028_ MuI._0372_ MuI._0614_ MuI._2789_ MuI._2791_ vssd1 vssd1 vccd1 vccd1 MuI._1874_
+ sky130_fd_sc_hd__and4_1
XFILLER_147_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ _02754_ _02797_ _05187_ _06518_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__and4_1
XFILLER_181_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08732__A _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07977__A1 _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07977__B2 _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ _00508_ _00509_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__nor2_1
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09547__B _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6587__B MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07016_ _05595_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__and3_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11525__A2 _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08967_ _01576_ _01577_ _01583_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__and3_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._706__B2 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07918_ _06522_ _00533_ _00535_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__or3_1
X_08898_ _01514_ _01515_ _06680_ _00085_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__and4bb_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4835__B MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07083__A _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__C _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07849_ _00236_ _00238_ _00239_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a21bo_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _03437_ _03439_ _03589_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__a211oi_4
XANTENNA__11036__C _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ _02146_ _02145_ _02144_ _02127_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o211a_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _03347_ _03345_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__or2b_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _02853_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10264__A2 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6041__A2 MuI._2889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _00292_ _06477_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nand2_1
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._105_ FuI._052_ FuI._060_ FuI._062_ FuI.a_operand\[11\] vssd1 vssd1 vccd1 vccd1
+ FuI._001_ sky130_fd_sc_hd__o31a_1
XANTENNA__13202__A2 _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _04085_ _04067_ _04069_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__nand3_1
X_12392_ _05130_ _05131_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__nor2_1
XFILLER_181_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11343_ _04110_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__xnor2_4
XFILLER_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ _04034_ _04036_ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__or3_1
XFILLER_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ _05822_ _05865_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12713__B2 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _02907_ _02908_ _02777_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__o21bai_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5304__A1 MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _05595_ _03454_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__or2b_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3660_ MuI._2605_ vssd1 vssd1 vccd1 vccd1 MuI._2616_ sky130_fd_sc_hd__clkbuf_4
XFILLER_208_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10087_ _02758_ _02759_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__nor2_2
XFILLER_75_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3591_ MuI._0592_ MuI._1285_ MuI._1846_ MuI._1824_ vssd1 vssd1 vccd1 vccd1 MuI._1857_
+ sky130_fd_sc_hd__a31o_1
XFILLER_63_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6018__A MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5330_ MuI._0969_ MuI._0970_ MuI._0971_ vssd1 vssd1 vccd1 vccd1 MuI._1106_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1204_ AuI._0263_ AuI._0408_ AuI._0288_ vssd1 vssd1 vccd1 vccd1 AuI._0409_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11543__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5261_ MuI._0912_ MuI._0920_ MuI._0919_ vssd1 vssd1 vccd1 vccd1 MuI._1030_ sky130_fd_sc_hd__a21bo_1
XAuI._1135_ AuI._0304_ AuI._0320_ AuI._0342_ vssd1 vssd1 vccd1 vccd1 AuI._0344_ sky130_fd_sc_hd__nor3b_2
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _03727_ _03728_ _03543_ _03547_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__o211ai_1
XMuI._4212_ MuI._3310_ MuI._3311_ vssd1 vssd1 vccd1 vccd1 MuI._3312_ sky130_fd_sc_hd__nor2_1
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5192_ MuI._0853_ MuI._0855_ MuI._0854_ vssd1 vssd1 vccd1 vccd1 MuI._0954_ sky130_fd_sc_hd__or3_1
XFILLER_31_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12728_ _03228_ _05820_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
XAuI._1066_ AuI._0228_ AuI._0238_ AuI._0175_ vssd1 vssd1 vccd1 vccd1 AuI._0277_ sky130_fd_sc_hd__mux2_1
XFILLER_203_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4480__B MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4143_ MuI._0361_ MuI._0614_ MuI._2330_ MuI._2830_ vssd1 vssd1 vccd1 vccd1 MuI._3243_
+ sky130_fd_sc_hd__and4_1
XFILLER_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ _05405_ _05412_ _05411_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._3808__C MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4074_ MuI._3160_ MuI._3171_ vssd1 vssd1 vccd1 vccd1 MuI._3174_ sky130_fd_sc_hd__nor2_1
XFILLER_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12401__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08552__A _01150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07168__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0919_ net131 net56 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0135_ sky130_fd_sc_hd__mux2_1
XANTENNA__09086__C _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4976_ MuI._1791_ MuI._0304_ MuI._0444_ MuI._1296_ vssd1 vssd1 vccd1 vccd1 MuI._0717_
+ sky130_fd_sc_hd__a22o_1
X_09870_ _02515_ _02511_ _02513_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__and3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6715_ MuI._2625_ MuI._2629_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2630_ sky130_fd_sc_hd__mux2_1
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3927_ MuI._2995_ MuI._3026_ vssd1 vssd1 vccd1 vccd1 MuI._3027_ sky130_fd_sc_hd__and2_1
XANTENNA__12180__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08821_ net111 _06581_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__nand2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__A _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6646_ MuI._1451_ MuI._1408_ vssd1 vssd1 vccd1 vccd1 MuI._2554_ sky130_fd_sc_hd__or2b_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3858_ MuI._2955_ MuI._2957_ vssd1 vssd1 vccd1 vccd1 MuI._2958_ sky130_fd_sc_hd__xnor2_1
X_08752_ _06593_ _04369_ _01354_ _01355_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__o2bb2a_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07703_ _00292_ _04111_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__nand2_1
XMuI._6577_ MuI._0680_ MuI._0713_ vssd1 vssd1 vccd1 vccd1 MuI._2478_ sky130_fd_sc_hd__nand2_1
XFILLER_66_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3789_ MuI.a_operand\[28\] MuI.a_operand\[27\] MuI.a_operand\[29\] MuI.a_operand\[30\]
+ vssd1 vssd1 vccd1 vccd1 MuI._2889_ sky130_fd_sc_hd__or4_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08683_ _01298_ _01299_ _01242_ _01300_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__and4bb_1
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5528_ MuI._1321_ MuI._1322_ MuI._1313_ MuI._1320_ vssd1 vssd1 vccd1 vccd1 MuI._1324_
+ sky130_fd_sc_hd__o211a_1
XFILLER_199_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07634_ _00121_ _00143_ _00250_ _00249_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__o211ai_2
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI.pe._408_ AuI.pe.significand\[5\] AuI.pe.significand\[4\] AuI.pe.significand\[6\]
+ AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 AuI.pe._375_ sky130_fd_sc_hd__or4_2
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5459_ MuI._2895_ MuI._0111_ vssd1 vssd1 vccd1 vccd1 MuI._1248_ sky130_fd_sc_hd__nand2_1
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07565_ _00173_ _00182_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__xor2_1
XANTENNA_MuI._4671__A MuI._1010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13432__A2 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _01913_ _01915_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10246__A2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07350__B _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _00109_ _00111_ _00110_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__o21ai_1
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ _01298_ _01299_ _01242_ _01300_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10992__A _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__A1 _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4585__A2 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09166_ _01775_ _01782_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a21oi_2
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08117_ _00237_ _00462_ _04778_ _04832_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__and4_1
XFILLER_147_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ net122 _00266_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nand2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07078__A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ _03820_ _03928_ _00516_ _00515_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a31o_1
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10706__B1 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _02665_ _02666_ _02676_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a21o_1
XFILLER_77_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06710__A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _02664_ _02663_ _02662_ _02659_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__o211ai_1
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3750__A MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0974__A1 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10232__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__D _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11961_ _04771_ _04775_ _04776_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand3_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__B1 _04843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _03473_ _03471_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and2b_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ _04700_ _04701_ _04551_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ _01146_ _00445_ _00550_ _01147_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a22oi_1
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10774_ _03493_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or2_1
XFILLER_198_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12513_ _02916_ _04929_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4731__D MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13493_ MuI.Underflow _02042_ _02151_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__and3_4
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13187__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12444_ _05203_ _05206_ _05204_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__o21ba_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _05181_ _05222_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__nor3_4
XFILLER_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__B _00708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _04026_ _04027_ _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__a211o_2
XFILLER_181_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6658__D MuI._2566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07419__C net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6020__B MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10126__B _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4830_ MuI._0552_ MuI._0555_ vssd1 vssd1 vccd1 vccd1 MuI._0556_ sky130_fd_sc_hd__and2b_1
XFILLER_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _04013_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__or2_1
XFILLER_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._690_ AuI.pe._211_ AuI.pe._385_ AuI.pe._208_ vssd1 vssd1 vccd1 vccd1 AuI.pe._238_
+ sky130_fd_sc_hd__or3_1
XFILLER_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4761_ MuI._0478_ MuI._0479_ MuI.b_operand\[11\] MuI._3223_ vssd1 vssd1 vccd1
+ vccd1 MuI._0480_ sky130_fd_sc_hd__and4bb_1
X_10208_ _02786_ _02772_ _02889_ _02784_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a31o_1
XFILLER_68_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12162__A2 _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output69_A net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09634__C _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ _03943_ _03944_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o211a_1
XMuI._6500_ MuI._1909_ MuI._1915_ MuI._1993_ vssd1 vssd1 vccd1 vccd1 MuI._2393_ sky130_fd_sc_hd__a21o_1
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3712_ MuI.b_operand\[19\] MuI._2811_ MuI._2773_ MuI._2786_ vssd1 vssd1 vccd1
+ vccd1 MuI._2812_ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3660__A MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4692_ MuI._0326_ MuI._0367_ vssd1 vssd1 vccd1 vccd1 MuI._0404_ sky130_fd_sc_hd__xor2_1
X_10139_ _03626_ _05788_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__or2_1
XFILLER_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6431_ MuI._2276_ MuI._2269_ vssd1 vssd1 vccd1 vccd1 MuI._2317_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3643_ MuI.a_operand\[13\] vssd1 vssd1 vccd1 vccd1 MuI._2429_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10499__D _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4906__D MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6362_ MuI._2239_ MuI._2240_ vssd1 vssd1 vccd1 vccd1 MuI._2241_ sky130_fd_sc_hd__or2_1
XFILLER_91_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3574_ MuI._1659_ MuI._1582_ vssd1 vssd1 vccd1 vccd1 MuI._1670_ sky130_fd_sc_hd__nor2_1
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5313_ MuI._1069_ MuI._1068_ vssd1 vssd1 vccd1 vccd1 MuI._1088_ sky130_fd_sc_hd__and2b_1
XANTENNA_MuI._6253__A2 MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__B _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6293_ MuI._2164_ MuI._1846_ vssd1 vssd1 vccd1 vccd1 MuI._2166_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13172__B _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4264__A1 MuI._1142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4264__B2 MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08266__B _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5244_ MuI._0938_ MuI._0937_ vssd1 vssd1 vccd1 vccd1 MuI._1012_ sky130_fd_sc_hd__and2b_1
XAuI._1118_ AuI._0326_ AuI._0327_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[2\]
+ sky130_fd_sc_hd__nor2_4
XFILLER_16_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07350_ _06544_ _05498_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__nand2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07601__D _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5175_ MuI._0934_ MuI._0935_ vssd1 vssd1 vccd1 vccd1 MuI._0936_ sky130_fd_sc_hd__nor2_1
XAuI._1049_ AuI._0254_ AuI._0260_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[0\]
+ sky130_fd_sc_hd__nor2_1
X_07281_ _06578_ _06579_ _06580_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__and4_1
XFILLER_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4126_ MuI._3224_ MuI._3225_ vssd1 vssd1 vccd1 vccd1 MuI._3226_ sky130_fd_sc_hd__nor2_1
XANTENNA__13178__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ _01635_ _01636_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a21o_1
XFILLER_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11728__A2 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4057_ MuI._3037_ MuI._3156_ vssd1 vssd1 vccd1 vccd1 MuI._3157_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09097__B _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10936__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09922_ _02575_ _02579_ _02580_ _02581_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a211o_1
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4959_ MuI._2841_ MuI._2352_ MuI._0591_ MuI._0593_ vssd1 vssd1 vccd1 vccd1 MuI._0698_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09853_ _02465_ _02464_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__and2b_1
XANTENNA__10061__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13347__B _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4666__A MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A2 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08804_ _01420_ _01421_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__xnor2_4
X_09784_ _02424_ _02432_ _02433_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nand3_1
XANTENNA__10052__A _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _05380_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13102__A1 _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6629_ MuI._1809_ MuI._1814_ MuI._1815_ vssd1 vssd1 vccd1 vccd1 MuI._2535_ sky130_fd_sc_hd__a21oi_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._753__A AuI.pe.significand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13102__B2 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _01348_ _01352_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3720__D MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09560__B _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08666_ _01281_ _01282_ _01283_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__o21bai_1
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08457__A _01071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _00233_ _00234_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__xor2_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _02420_ _06513_ _06602_ _06604_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__and4_1
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11416__A1 _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07548_ _00161_ _00165_ vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__nor2_1
XFILLER_167_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09085__A2 _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07479_ _00095_ _00096_ _04509_ _00035_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__and4_1
XFILLER_210_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08832__A2 _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13169__A1 _04678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ _01729_ _01730_ _01731_ _01711_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__o22a_1
XANTENNA__11611__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ _03007_ _03015_ _03014_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06705__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12426__B _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12916__A1 _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3745__A MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _01679_ _01766_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12916__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11330__B _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1436__A2 AuI._0519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ _04989_ _04990_ _04904_ _04862_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__o211a_2
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08342__D net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3518__B1 MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11111_ _03738_ _03739_ _03816_ _03817_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__nor4b_1
XFILLER_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _04915_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12442__A _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4730__A2 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11042_ _06680_ _00382_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3480__A MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input20_A a_operand[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10897__A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ _03550_ _03615_ _05660_ _05713_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__and4_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13273__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _04604_ _04610_ _04757_ _04758_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a211o_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ _03152_ _06666_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nand2_1
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10826_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__nor2_1
XFILLER_158_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11958__A2 _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4461__D MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _03280_ _03283_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__nor2_1
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1675__A2 AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _00955_ _00956_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nor2_1
X_10688_ _03404_ _03405_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__and3_1
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12427_ _05276_ _05277_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__or3_1
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5931_ MuI._1717_ MuI._1754_ vssd1 vssd1 vccd1 vccd1 MuI._1767_ sky130_fd_sc_hd__or2b_1
XFILLER_127_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _05203_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__nor2_1
XFILLER_153_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._811_ AuI.pe._095_ AuI.pe._370_ AuI.pe._349_ AuI.pe._336_ AuI.pe._337_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._350_ sky130_fd_sc_hd__o221a_1
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5862_ MuI._2790_ MuI._0168_ MuI._0683_ MuI._0684_ vssd1 vssd1 vccd1 vccd1 MuI._1691_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _00095_ _00096_ _05241_ _05305_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__and4_2
XFILLER_206_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12289_ _04991_ _04993_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__nor2_1
XFILLER_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._742_ AuI.pe._145_ AuI.pe._388_ AuI.pe._286_ vssd1 vssd1 vccd1 vccd1 AuI.pe._287_
+ sky130_fd_sc_hd__and3_1
XMuI._4813_ MuI._0403_ MuI._0404_ vssd1 vssd1 vccd1 vccd1 MuI._0538_ sky130_fd_sc_hd__xor2_1
XMuI._5793_ MuI._2429_ MuI._3306_ MuI._2881_ MuI._2660_ vssd1 vssd1 vccd1 vccd1 MuI._1616_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1667_ AuI.operand_a\[28\] AuI._0604_ AuI._0692_ AuI.operand_a\[29\] AuI._0258_
+ vssd1 vssd1 vccd1 vccd1 AuI._0019_ sky130_fd_sc_hd__a311o_1
XAuI.pe._673_ AuI.pe._170_ AuI.pe._050_ AuI.pe._220_ AuI.pe._221_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._222_ sky130_fd_sc_hd__a211o_1
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4744_ MuI._0458_ MuI._0461_ vssd1 vssd1 vccd1 vccd1 MuI._0462_ sky130_fd_sc_hd__nor2_1
XFILLER_95_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ _03809_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__clkbuf_4
XAuI._1598_ AuI._0259_ AuI._0768_ AuI._0770_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[13\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4675_ MuI._0380_ MuI._0384_ vssd1 vssd1 vccd1 vccd1 MuI._0386_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06781_ _03067_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__and3_1
XANTENNA__13096__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5682__B1 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6414_ MuI._2153_ MuI._2298_ vssd1 vssd1 vccd1 vccd1 MuI._2299_ sky130_fd_sc_hd__nor2_1
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3626_ MuI._1538_ MuI._1549_ vssd1 vssd1 vccd1 vccd1 MuI._2242_ sky130_fd_sc_hd__and2_1
X_08520_ _01102_ _01098_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__and2b_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6345_ MuI._2221_ MuI._2222_ vssd1 vssd1 vccd1 vccd1 MuI._2223_ sky130_fd_sc_hd__xor2_1
XMuI._3557_ MuI._1472_ vssd1 vssd1 vccd1 vccd1 MuI._1483_ sky130_fd_sc_hd__clkbuf_4
X_08451_ _00883_ _00885_ _00884_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__o21ai_1
XFILLER_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11415__B _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5434__B1 MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07612__C _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5748__C MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13399__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07402_ _00018_ _00016_ _00017_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__nand3_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6276_ MuI._2054_ MuI._2050_ vssd1 vssd1 vccd1 vccd1 MuI._2147_ sky130_fd_sc_hd__and2b_1
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3549__B MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3488_ MuI._0680_ MuI._0713_ vssd1 vssd1 vccd1 vccd1 MuI._0724_ sky130_fd_sc_hd__xnor2_1
X_08382_ _00996_ _00998_ _00997_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a21o_1
XFILLER_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5227_ MuI._0896_ MuI._0902_ vssd1 vssd1 vccd1 vccd1 MuI._0993_ sky130_fd_sc_hd__or2b_1
X_07333_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__nor2_1
XANTENNA__12071__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5158_ MuI._0914_ MuI._0915_ MuI._0916_ vssd1 vssd1 vccd1 vccd1 MuI._0917_ sky130_fd_sc_hd__or3_1
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5764__B MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _06564_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4109_ MuI._3206_ MuI._3208_ vssd1 vssd1 vccd1 vccd1 MuI._3209_ sky130_fd_sc_hd__and2_1
X_09003_ _01436_ _01618_ _01619_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nand4b_1
XANTENNA__13034__A1_N _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5089_ MuI._0806_ MuI._0814_ MuI._0827_ vssd1 vssd1 vccd1 vccd1 MuI._0841_ sky130_fd_sc_hd__and3_1
X_07195_ _06494_ _06495_ net21 _06461_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__and4_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._143__149 vssd1 vssd1 vccd1 vccd1 FuI._143__149/HI net149 sky130_fd_sc_hd__conb_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6162__A1 MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6162__B2 MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09905_ _02530_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__and2_1
XFILLER_86_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09836_ _02477_ _02479_ _02438_ _02480_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a211o_1
XANTENNA__11309__C _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09767_ _02248_ _00287_ _02361_ _02360_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
X_06979_ _05198_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__clkbuf_4
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09290__B _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _01333_ _01335_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__nor2_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _02166_ _02218_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__and2_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__B1 _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07091__A _04929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08649_ _01262_ _01264_ _01266_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__or3_2
XFILLER_203_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6116__A MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ _04449_ _04452_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__nand3_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _03319_ _03321_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a21o_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12062__B2 _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ _04373_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__xor2_1
XFILLER_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13330_ _06239_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__nor2_1
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ _02539_ _05649_ _03246_ _03248_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nand4_1
XFILLER_183_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5674__B MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3475__A MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _03669_ _05842_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__nand2_1
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _02994_ _02996_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__nor2_1
XFILLER_6_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _05045_ _05046_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _02837_ _06097_ _02713_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__a21oi_1
XFILLER_151_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input68_A b_operand[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__B2 _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _04970_ _04971_ _04839_ _04844_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__o211a_1
XFILLER_151_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1521_ AuI._0701_ AuI._0612_ AuI._0703_ AuI._0705_ vssd1 vssd1 vccd1 vccd1 AuI._0706_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07266__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__clkinv_2
XANTENNA__08800__D _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__C _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _03768_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__and2b_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1452_ AuI._0462_ AuI._0467_ vssd1 vssd1 vccd1 vccd1 AuI._0638_ sky130_fd_sc_hd__xor2_2
XFILLER_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4467__A1 MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1383_ AuI._0559_ AuI._0564_ vssd1 vssd1 vccd1 vccd1 AuI._0574_ sky130_fd_sc_hd__nor2_1
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4467__B2 MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6725__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4460_ MuI.a_operand\[20\] MuI.b_operand\[1\] MuI.b_operand\[0\] MuI.a_operand\[21\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0149_ sky130_fd_sc_hd__a22o_1
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._521__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__A _00810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _03454_ _05831_ _05895_ _03389_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a22oi_1
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4391_ MuI._0049_ MuI._0050_ vssd1 vssd1 vccd1 vccd1 MuI._0074_ sky130_fd_sc_hd__and2b_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _04721_ _04740_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nand3_1
XFILLER_61_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6130_ MuI._1904_ MuI._1906_ vssd1 vssd1 vccd1 vccd1 MuI._1986_ sky130_fd_sc_hd__or2b_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11858_ _03013_ _05660_ _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__nand4_1
XMuI._6061_ MuI._3036_ MuI._3035_ vssd1 vssd1 vccd1 vccd1 MuI._1910_ sky130_fd_sc_hd__and2b_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _03399_ _03408_ _03407_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__a21o_1
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11789_ _04420_ _04422_ _04591_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__o211ai_4
XMuI._5012_ MuI._0686_ MuI._0688_ vssd1 vssd1 vccd1 vccd1 MuI._0756_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5584__B MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0856__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5195__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ _06372_ _06373_ _02700_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__o21bai_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__A2 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09656__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5914_ MuI._1741_ MuI._1742_ MuI._1746_ MuI._1748_ vssd1 vssd1 vccd1 vccd1 MuI._1749_
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13305__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5845_ MuI._0696_ MuI._1672_ vssd1 vssd1 vccd1 vccd1 MuI._1673_ sky130_fd_sc_hd__nor2_1
XANTENNA__07176__A _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ _00051_ _00568_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__nor2_1
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._725_ AuI.pe._386_ AuI.pe._238_ AuI.pe.significand\[20\] vssd1 vssd1 vccd1
+ vccd1 AuI.pe._271_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06902_ _04369_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_MuI._5105__A MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5776_ MuI._1518_ MuI._1536_ MuI._1537_ vssd1 vssd1 vccd1 vccd1 MuI._1597_ sky130_fd_sc_hd__nand3_1
X_07882_ _00343_ _00357_ _00356_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__o21ba_1
XFILLER_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._656_ AuI.pe._084_ AuI.pe._112_ AuI.pe._199_ AuI.pe._205_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._206_ sky130_fd_sc_hd__a211o_1
XMuI._4727_ MuI._0309_ MuI._0442_ vssd1 vssd1 vccd1 vccd1 MuI._0443_ sky130_fd_sc_hd__or2_1
XANTENNA__08805__B_N _01422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06833_ _03626_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__and3_1
X_09621_ _02253_ _02256_ _02208_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__o211ai_2
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._587_ AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 AuI.pe._142_ sky130_fd_sc_hd__buf_2
XANTENNA__08719__B _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4658_ MuI._0364_ MuI._0366_ vssd1 vssd1 vccd1 vccd1 MuI._0367_ sky130_fd_sc_hd__xnor2_1
X_09552_ _02082_ _02084_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10330__A _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06764_ net43 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__buf_4
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09541__D _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3609_ MuI.a_operand\[17\] vssd1 vssd1 vccd1 vccd1 MuI._2055_ sky130_fd_sc_hd__clkbuf_4
X_08503_ _00848_ _00847_ _00846_ _00835_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__o211a_1
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4589_ MuI._0219_ MuI._0289_ MuI._0290_ vssd1 vssd1 vccd1 vccd1 MuI._0291_ sky130_fd_sc_hd__or3_1
XANTENNA__11095__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _01975_ _01974_ _01973_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__o21ai_1
X_06695_ _02140_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__buf_2
XANTENNA__07342__C net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6328_ MuI._2173_ MuI._2174_ MuI._2177_ MuI._2203_ MuI._2182_ vssd1 vssd1 vccd1
+ vccd1 MuI._2204_ sky130_fd_sc_hd__o32a_1
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08434_ _00835_ _00845_ _00844_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1386__S AuI._0126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6259_ MuI._0328_ MuI._2894_ MuI._2550_ MuI._2517_ vssd1 vssd1 vccd1 vccd1 MuI._2128_
+ sky130_fd_sc_hd__and4_1
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _00971_ _00976_ _00972_ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI._1639__A2 AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08454__B _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _06524_ _06530_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__or2b_1
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08799__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08296_ _03346_ _03982_ _00912_ _00913_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__a31o_1
XANTENNA__09269__C net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08173__C net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ net109 vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__buf_4
XFILLER_164_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._579__A2 AuI.pe._026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ net110 vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__buf_4
XFILLER_180_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10358__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10358__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09285__B _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06702__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09716__D _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3742__B MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5894__B1 MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _02469_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__or2_1
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07533__B _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _05624_ _05626_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2b_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05635_ _05636_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__xnor2_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11712_ _04371_ _04500_ _04508_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a21oi_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__A2 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _05561_ _05562_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__and2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _04433_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__xor2_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or2_1
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10597__A1 _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 a_operand[20] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_6
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10597__B2 _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 a_operand[30] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
XFILLER_183_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 b_operand[11] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_4
X_10525_ _03230_ _03227_ _03229_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__nand3_1
X_13313_ _06194_ _06166_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__or2b_1
XAuI._0952_ AuI._0163_ vssd1 vssd1 vccd1 vccd1 AuI._0164_ sky130_fd_sc_hd__clkbuf_2
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _02645_ _06089_ _02687_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__a21o_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10456_ _03155_ _03156_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__xnor2_4
XAuI._0883_ AuI._0035_ AuI._0095_ AuI._0102_ vssd1 vssd1 vccd1 vccd1 AuI._0103_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11546__B1 _02719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3960_ MuI._3039_ MuI._3053_ MuI._3054_ MuI._3059_ vssd1 vssd1 vccd1 vccd1 MuI._3060_
+ sky130_fd_sc_hd__or4b_1
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ _06075_ _06077_ _06080_ _02841_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a31o_1
X_10387_ net108 _05756_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__and2_1
X_12126_ net61 _04854_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__nand2_1
XMuI._3891_ MuI._2913_ MuI._2922_ vssd1 vssd1 vccd1 vccd1 MuI._2991_ sky130_fd_sc_hd__and2_1
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13299__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07427__C _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5630_ MuI._1426_ MuI._1435_ vssd1 vssd1 vccd1 vccd1 MuI._1436_ sky130_fd_sc_hd__nor2_1
XAuI._1504_ AuI._0688_ AuI._0689_ vssd1 vssd1 vccd1 vccd1 AuI._0690_ sky130_fd_sc_hd__nor2_1
X_12057_ _02575_ _02579_ _03315_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__o21ai_1
XFILLER_96_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11849__A1 _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._510_ AuI.pe.significand\[6\] AuI.pe._065_ vssd1 vssd1 vccd1 vccd1 AuI.pe._070_
+ sky130_fd_sc_hd__or2_2
XANTENNA__12630__A _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__D _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5561_ MuI._1343_ MuI._1358_ MuI._1359_ vssd1 vssd1 vccd1 vccd1 MuI._1360_ sky130_fd_sc_hd__o21ba_1
X_11008_ _03748_ _03749_ _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a21o_1
XAuI._1435_ AuI._0504_ AuI._0506_ vssd1 vssd1 vccd1 vccd1 AuI._0621_ sky130_fd_sc_hd__and2_1
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._441_ AuI.pe.significand\[8\] vssd1 vssd1 vccd1 vccd1 AuI.pe._008_ sky130_fd_sc_hd__inv_2
XANTENNA__10521__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4512_ MuI._0183_ MuI._0204_ MuI._0205_ vssd1 vssd1 vccd1 vccd1 MuI._0206_ sky130_fd_sc_hd__a21o_1
XANTENNA__10521__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1030__A3 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11246__A _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5492_ MuI._1276_ MuI._1282_ MuI._1283_ vssd1 vssd1 vccd1 vccd1 MuI._1284_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._5101__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07443__B _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5579__B MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1366_ AuI._0539_ AuI._0540_ AuI._0546_ AuI._0557_ vssd1 vssd1 vccd1 vccd1 AuI._0559_
+ sky130_fd_sc_hd__nand4_2
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4443_ MuI._0128_ MuI._0129_ vssd1 vssd1 vccd1 vccd1 MuI._0131_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _03306_ _02809_ _05849_ _03239_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a2bb2o_1
XAuI._1297_ AuI._0484_ AuI._0485_ AuI._0494_ AuI._0495_ vssd1 vssd1 vccd1 vccd1 AuI._0496_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4374_ MuI._0052_ MuI._0053_ MuI._0055_ vssd1 vssd1 vccd1 vccd1 MuI._0056_ sky130_fd_sc_hd__o21ba_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6113_ MuI._1887_ MuI._1888_ vssd1 vssd1 vccd1 vccd1 MuI._1968_ sky130_fd_sc_hd__and2_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6044_ MuI._3129_ MuI._3131_ vssd1 vssd1 vccd1 vccd1 MuI._1892_ sky130_fd_sc_hd__nand2_1
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _00419_ _00428_ _00766_ _00767_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__a211o_1
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ _06056_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__clkbuf_2
XFILLER_147_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _00696_ _00697_ _00693_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__a21o_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ _05767_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__clkbuf_4
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11001__A2 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07618__B _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6877_ MuI._2735_ MuI._2776_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[29\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_103_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _01597_ _01592_ _01593_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__nand3_1
XANTENNA__10044__B _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5828_ MuI._1584_ MuI._1586_ MuI._1585_ vssd1 vssd1 vccd1 vccd1 MuI._1654_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1006__A0 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _06587_ _00551_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__nor2_1
XAuI.pe._708_ AuI.pe._074_ AuI.pe._241_ AuI.pe._243_ AuI.pe._254_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[19\] sky130_fd_sc_hd__o22a_1
XFILLER_111_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5759_ MuI._1575_ MuI._1576_ MuI._1577_ vssd1 vssd1 vccd1 vccd1 MuI._1578_ sky130_fd_sc_hd__nand3b_1
X_07865_ _00249_ _00252_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__nand2_1
XAuI.pe._639_ AuI.pe._120_ AuI.pe._025_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._190_
+ sky130_fd_sc_hd__a21o_1
X_09604_ _02221_ _02220_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__and2b_1
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10060__A _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _03443_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__clkbuf_8
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07796_ net68 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__buf_6
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08168__C _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _02164_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__nor2_1
X_06747_ net39 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__buf_6
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__and2_1
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08417_ _01027_ _01034_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__nand2_1
XFILLER_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09397_ _02012_ _02013_ _02003_ _02008_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a211o_1
XANTENNA_MuI._4603__B2 MuI._2939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._121_ FuI._023_ FuI._054_ FuI._058_ FuI.a_operand\[17\] vssd1 vssd1 vccd1 vccd1
+ FuI._031_ sky130_fd_sc_hd__o31a_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12568__A2 _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _06500_ _06517_ _06518_ _06501_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._3957__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFuI._149__155 vssd1 vssd1 vccd1 vccd1 FuI._149__155/HI net155 sky130_fd_sc_hd__conb_1
XANTENNA__10219__B _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _00892_ _00893_ _00896_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__or3_1
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11041__D net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13310__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _02998_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__xnor2_2
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11290_ _03922_ _03925_ _03923_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__o21bai_1
XANTENNA__06713__A _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__D _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3753__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__buf_4
XFILLER_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09446__D net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3472__B MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _02850_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__inv_2
XFILLER_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10889__B _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07544__A _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4584__A MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__A2 _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1220_ AuI._0210_ AuI._0423_ AuI._0389_ vssd1 vssd1 vccd1 vccd1 AuI._0424_ sky130_fd_sc_hd__mux2_1
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1151_ AuI._0344_ AuI._0358_ vssd1 vssd1 vccd1 vccd1 AuI._0359_ sky130_fd_sc_hd__or2_1
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12256__A1 _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ _03346_ _05842_ _05690_ _05691_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12256__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _03486_ _05585_ _05616_ _05617_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand4_1
XAuI._1082_ AuI._0185_ AuI._0292_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0293_ sky130_fd_sc_hd__mux2_1
XFILLER_203_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08375__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08806__C _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _05543_ _05544_ _05455_ _05458_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a211o_1
XFILLER_203_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4750__C MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4090_ MuI.b_operand\[6\] vssd1 vssd1 vccd1 vccd1 MuI._3190_ sky130_fd_sc_hd__clkbuf_4
X_11626_ _04398_ _04399_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__a21o_1
XFILLER_156_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11557_ _02771_ _04175_ _02772_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12625__A _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A2 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10508_ _03195_ _03197_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a21o_1
XAuI._0935_ AuI._0143_ AuI._0146_ AuI._0100_ vssd1 vssd1 vccd1 vccd1 AuI._0147_ sky130_fd_sc_hd__a21o_1
XANTENNA__07719__A _06455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output99_A net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _04267_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__xnor2_4
XANTENNA_MuI._4759__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6800_ MuI._2630_ MuI._2680_ MuI._2632_ vssd1 vssd1 vccd1 vccd1 MuI._2723_ sky130_fd_sc_hd__o21bai_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12344__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3663__A MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4992_ MuI._0733_ vssd1 vssd1 vccd1 vccd1 MuI._0734_ sky130_fd_sc_hd__inv_2
X_10439_ _02977_ _03000_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__a21boi_2
X_13227_ _06029_ _06032_ _06133_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nand3_1
XAuI._0866_ AuI._0056_ AuI._0066_ AuI._0077_ AuI._0085_ vssd1 vssd1 vccd1 vccd1 AuI._0086_
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4478__B MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6731_ MuI._2640_ MuI._2646_ MuI._2487_ vssd1 vssd1 vccd1 vccd1 MuI._2647_ sky130_fd_sc_hd__mux2_1
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12192__B1 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3943_ MuI._3040_ MuI._3041_ MuI._3042_ vssd1 vssd1 vccd1 vccd1 MuI._3043_ sky130_fd_sc_hd__or3_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13158_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__nor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6662_ MuI._2509_ MuI._2570_ MuI._2485_ vssd1 vssd1 vccd1 vccd1 MuI._2571_ sky130_fd_sc_hd__mux2_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3874_ MuI._0768_ MuI._1010_ MuI._2844_ MuI._2838_ vssd1 vssd1 vccd1 vccd1 MuI._2974_
+ sky130_fd_sc_hd__and4_1
X_12109_ _04935_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ _05918_ _05922_ _05915_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__o21a_1
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._5613_ MuI._1415_ MuI._1416_ MuI._3269_ MuI._0420_ vssd1 vssd1 vccd1 vccd1 MuI._1418_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07454__A net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6593_ MuI._0273_ MuI._2493_ MuI._2494_ vssd1 vssd1 vccd1 vccd1 MuI._2496_ sky130_fd_sc_hd__a21o_1
XANTENNA_AuI._1502__B AuI._0586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4494__A MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5544_ MuI._2876_ MuI._0321_ MuI._1335_ MuI._1339_ vssd1 vssd1 vccd1 vccd1 MuI._1342_
+ sky130_fd_sc_hd__a211oi_1
XAuI._1418_ AuI.operand_a\[30\] AuI.operand_a\[28\] AuI.operand_a\[29\] AuI._0604_
+ vssd1 vssd1 vccd1 vccd1 AuI._0605_ sky130_fd_sc_hd__and4_1
X_07650_ _03217_ _03271_ _00267_ _04294_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__and4_1
XFILLER_26_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._424_ AuI.pe._382_ AuI.pe._384_ AuI.pe._387_ AuI.pe._390_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._391_ sky130_fd_sc_hd__and4_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._479__A1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5475_ MuI._2874_ MuI._2876_ MuI._0315_ MuI.a_operand\[0\] vssd1 vssd1 vccd1
+ vccd1 MuI._1266_ sky130_fd_sc_hd__and4_1
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1349_ AuI._0538_ AuI._0541_ AuI._0542_ vssd1 vssd1 vccd1 vccd1 AuI._0544_ sky130_fd_sc_hd__a21o_1
XFILLER_92_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _06601_ _06584_ _05112_ _06606_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a22o_1
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4519__A1_N MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4426_ MuI._0111_ vssd1 vssd1 vccd1 vccd1 MuI._0112_ sky130_fd_sc_hd__clkbuf_4
X_09320_ _01822_ _01821_ _01814_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a21o_1
XANTENNA__11704__A _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B _00518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4357_ MuI._0035_ MuI._0036_ vssd1 vssd1 vccd1 vccd1 MuI._0037_ sky130_fd_sc_hd__xor2_2
X_09251_ _01655_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__clkinv_2
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10608__A_N _03993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ _00162_ _06518_ _00412_ _00164_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__a22oi_2
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4288_ MuI._3385_ MuI._3383_ vssd1 vssd1 vccd1 vccd1 MuI._3388_ sky130_fd_sc_hd__xnor2_1
X_09182_ _02970_ _03895_ _03982_ _02916_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a22oi_1
XFILLER_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6027_ MuI._0625_ MuI._2789_ MuI._2791_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._1873_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08133_ _06601_ _05187_ _06568_ _06606_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__a22oi_1
XFILLER_174_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout120_A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08732__B _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07977__A2 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _00680_ _00681_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07015_ _05585_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08966_ _01576_ _01577_ _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07917_ _02528_ _00534_ _06514_ _06521_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12486__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ _06622_ _00035_ _04638_ _00414_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22oi_1
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12420__D _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _00463_ _00464_ _00461_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__D _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _06516_ _05498_ _05563_ _06520_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a22o_1
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _02127_ _02144_ _02145_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a211oi_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _03379_ _03415_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a21o_1
XANTENNA__06708__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11333__B _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09449_ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__inv_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6041__A3 MuI._2890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _05312_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nor2_1
XFuI._104_ FuI._037_ FuI._061_ FuI._056_ vssd1 vssd1 vccd1 vccd1 FuI._062_ sky130_fd_sc_hd__and3b_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08923__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11411_ _04052_ _04053_ _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__or4_2
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12391_ _05238_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__or2_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10421__B1 _03119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ _00502_ _04467_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__nand2_1
XFILLER_180_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11273_ _02712_ _03247_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__nand2_1
XANTENNA_input50_A b_operand[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4760__B1 MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12713__A2 _03974_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10224_ _02777_ _02778_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__or2_2
X_13012_ _05904_ _05905_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and2_1
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5304__A2 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _02831_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__nor2_2
XFILLER_95_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ _02388_ _04262_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__and2b_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3590_ MuI._1824_ MuI._1835_ vssd1 vssd1 vccd1 vccd1 MuI._1846_ sky130_fd_sc_hd__nor2_1
XANTENNA__10156__B_N _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__C1 _04481_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6018__B MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1203_ AuI._0273_ AuI._0290_ AuI._0291_ AuI._0293_ AuI._0274_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0408_ sky130_fd_sc_hd__mux4_1
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5260_ MuI._1027_ MuI._1028_ vssd1 vssd1 vccd1 vccd1 MuI._1029_ sky130_fd_sc_hd__nor2_1
XAuI._1134_ AuI._0304_ AuI._0320_ AuI._0342_ vssd1 vssd1 vccd1 vccd1 AuI._0343_ sky130_fd_sc_hd__o21bai_1
XFILLER_204_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4211_ MuI._1021_ MuI._2895_ vssd1 vssd1 vccd1 vccd1 MuI._3311_ sky130_fd_sc_hd__nand2_1
XANTENNA__11819__A1_N _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ _03543_ _03547_ _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a211o_1
XMuI._5191_ MuI._0928_ MuI._0929_ MuI._0950_ MuI._0951_ vssd1 vssd1 vccd1 vccd1 MuI._0953_
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA_MuI._3658__A MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12727_ _05551_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__inv_2
XAuI._1065_ AuI._0233_ vssd1 vssd1 vccd1 vccd1 AuI._0276_ sky130_fd_sc_hd__buf_2
XFILLER_203_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4142_ MuI._0614_ MuI._2330_ MuI._2830_ MuI._0361_ vssd1 vssd1 vccd1 vccd1 MuI._3242_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4480__C MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12658_ _05525_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__xor2_1
XANTENNA__08833__A _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3808__D MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4073_ MuI._2835_ MuI._2953_ vssd1 vssd1 vccd1 vccd1 MuI._3173_ sky130_fd_sc_hd__xor2_1
X_11609_ _04395_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a21o_1
XFILLER_191_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12401__B2 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _05444_ _05451_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nand3_2
XFILLER_184_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12952__A2 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0918_ AuI._0134_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[26\] sky130_fd_sc_hd__clkbuf_2
XANTENNA_AuI._1209__B1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09086__D _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4975_ MuI._0624_ MuI._0714_ MuI._0715_ vssd1 vssd1 vccd1 vccd1 MuI._0716_ sky130_fd_sc_hd__or3_1
XFILLER_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._0849_ AuI._0067_ net11 AuI._0068_ net10 vssd1 vssd1 vccd1 vccd1 AuI._0069_ sky130_fd_sc_hd__a22o_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__B1 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3926_ MuI._3011_ MuI._3025_ vssd1 vssd1 vccd1 vccd1 MuI._3026_ sky130_fd_sc_hd__xnor2_1
XMuI._6714_ MuI._2306_ MuI._2628_ vssd1 vssd1 vccd1 vccd1 MuI._2629_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08820_ _02096_ _02194_ net14 net15 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__and4_1
XFILLER_98_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__A _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6645_ MuI._2547_ MuI._2552_ vssd1 vssd1 vccd1 vccd1 MuI._2553_ sky130_fd_sc_hd__nor2_1
XFILLER_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3857_ MuI._2956_ MuI._2949_ vssd1 vssd1 vccd1 vccd1 MuI._2957_ sky130_fd_sc_hd__nor2_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _01366_ _01368_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__nor2_1
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6576_ MuI._2476_ vssd1 vssd1 vccd1 vccd1 MuI._2477_ sky130_fd_sc_hd__inv_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07702_ _00073_ _00076_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__nor2_1
XMuI._3788_ MuI._2883_ MuI._2887_ vssd1 vssd1 vccd1 vccd1 MuI._2888_ sky130_fd_sc_hd__nor2_1
XFILLER_39_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08682_ _01228_ _01241_ _01236_ _01240_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__a211o_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07344__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5527_ MuI._1313_ MuI._1320_ MuI._1321_ MuI._1322_ vssd1 vssd1 vccd1 vccd1 MuI._1323_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07912__A _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _00249_ _00250_ _00143_ _00121_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__a211o_1
XFILLER_199_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._407_ AuI.pe.significand\[8\] AuI.pe._372_ AuI.pe._373_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._374_ sky130_fd_sc_hd__or3_2
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5458_ MuI._1245_ MuI._1246_ vssd1 vssd1 vccd1 vccd1 MuI._1247_ sky130_fd_sc_hd__nor2_1
XANTENNA__11434__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _00180_ _00181_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__and2b_1
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4671__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4409_ MuI._3353_ MuI._3354_ vssd1 vssd1 vccd1 vccd1 MuI._0093_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09303_ _01919_ _01920_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__nand2_1
XMuI._5389_ MuI._1121_ MuI._1167_ MuI._1170_ vssd1 vssd1 vccd1 vccd1 MuI._1171_ sky130_fd_sc_hd__o21a_1
XANTENNA__10246__A3 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07495_ _06629_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__o21bai_1
XFILLER_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09839__A _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _01631_ _01632_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__and4bb_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5231__A1 MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10580__A_N _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5231__B2 MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ _01720_ _01722_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13196__A2 _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08116_ _03099_ _04778_ _06603_ _03056_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__a22oi_4
XFILLER_175_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09096_ net68 net38 net123 net34 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__and4_1
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4399__A MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08047_ _06458_ _00663_ _00664_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a21boi_2
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3545__A1 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10706__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10706__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5298__A1 MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__B_N _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06710__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _02659_ _02662_ _02663_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a211o_2
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__A2_N _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08949_ _01565_ _01564_ _01532_ _01508_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07525__C _00141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11960_ _04774_ _04773_ _04772_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__a21bo_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._753__C_N AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11131__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11131__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08532__C1 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _03558_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__xnor2_2
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4862__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _04551_ _04700_ _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or3_2
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10842_ _03568_ _03569_ _03570_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__a21o_1
XFILLER_60_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3478__A MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _03494_ _03318_ _03496_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__a211o_1
XFILLER_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12512_ _02621_ _05368_ _02619_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__and3_1
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5222__A1 MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ _04161_ _06385_ _06386_ _06403_ _06407_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__a311o_4
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _05294_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09468__B _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12395__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _05219_ _05221_ _05182_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o21a_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ _04052_ _04053_ _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__nor4_2
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4102__A MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__B1 _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07419__D _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11256_ _04014_ _04016_ _04019_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__or3_1
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06901__A _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3941__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4760_ MuI._2854_ MuI._0477_ MuI._2790_ MuI._2836_ vssd1 vssd1 vccd1 vccd1 MuI._0479_
+ sky130_fd_sc_hd__a22oi_1
X_10207_ _02879_ _02886_ _02757_ _02887_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a311o_1
X_11187_ _03907_ _03908_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a211oi_2
XFILLER_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3711_ MuI.b_operand\[18\] vssd1 vssd1 vccd1 vccd1 MuI._2811_ sky130_fd_sc_hd__clkbuf_2
XFILLER_121_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09634__D _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__A2_N _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4691_ MuI._0401_ MuI._0402_ vssd1 vssd1 vccd1 vccd1 MuI._0403_ sky130_fd_sc_hd__xor2_1
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _03615_ _05777_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__nand2_2
XFILLER_95_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6430_ MuI._2313_ MuI._2314_ MuI._1939_ MuI._2311_ vssd1 vssd1 vccd1 vccd1 MuI._2316_
+ sky130_fd_sc_hd__o211a_1
XMuI._3642_ MuI._2330_ MuI._0460_ MuI._2396_ MuI._2407_ MuI._2385_ vssd1 vssd1 vccd1
+ vccd1 MuI._2418_ sky130_fd_sc_hd__a32o_1
XFILLER_10_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10069_ _02706_ _02129_ _02064_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__and3b_1
XFILLER_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6238__B1 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6361_ MuI._2237_ MuI._2238_ MuI._2194_ MuI._2199_ vssd1 vssd1 vccd1 vccd1 MuI._2240_
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3573_ MuI._1076_ vssd1 vssd1 vccd1 vccd1 MuI._1659_ sky130_fd_sc_hd__inv_2
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5312_ MuI._0964_ MuI._0961_ MuI._0963_ vssd1 vssd1 vccd1 vccd1 MuI._1086_ sky130_fd_sc_hd__a21o_1
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6292_ MuI._0581_ MuI._1285_ vssd1 vssd1 vccd1 vccd1 MuI._2164_ sky130_fd_sc_hd__nand2_1
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4264__A2 MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4491__B MuI._0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5243_ MuI._0993_ MuI._0994_ MuI._1008_ vssd1 vssd1 vccd1 vccd1 MuI._1011_ sky130_fd_sc_hd__nand3_1
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1117_ AuI._0324_ AuI._0325_ vssd1 vssd1 vccd1 vccd1 AuI._0327_ sky130_fd_sc_hd__nor2_1
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5174_ MuI._2838_ MuI._0100_ MuI._0228_ MuI._2844_ vssd1 vssd1 vccd1 vccd1 MuI._0935_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ net13 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__clkbuf_4
XAuI._1048_ AuI._0259_ AuI._0252_ AuI._0140_ vssd1 vssd1 vccd1 vccd1 AuI._0260_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A _00934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4125_ MuI._1802_ MuI._2773_ MuI._2786_ MuI._2550_ vssd1 vssd1 vccd1 vccd1 MuI._3225_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_176_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13178__A2 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4056_ MuI._3154_ MuI._3155_ vssd1 vssd1 vccd1 vccd1 MuI._3156_ sky130_fd_sc_hd__nor2_1
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07179__A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _02484_ _02578_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__nor2_1
XANTENNA__06811__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4958_ MuI._0694_ MuI._0696_ vssd1 vssd1 vccd1 vccd1 MuI._0697_ sky130_fd_sc_hd__nor2_1
XANTENNA__11429__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _02505_ _02506_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__or2b_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3909_ MuI._2928_ MuI._2933_ vssd1 vssd1 vccd1 vccd1 MuI._3009_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._4666__B MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _01390_ _01389_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__and2b_1
XMuI._4889_ MuI._0432_ MuI._0619_ MuI._0620_ vssd1 vssd1 vccd1 vccd1 MuI._0621_ sky130_fd_sc_hd__or3_1
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _02407_ _02408_ _02423_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a21o_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _05370_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__buf_4
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6628_ MuI._2519_ MuI._2520_ MuI._2522_ MuI._2525_ MuI._2533_ vssd1 vssd1 vccd1
+ vccd1 MuI._2534_ sky130_fd_sc_hd__a2111o_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._753__B AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__A2 _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _01349_ _01350_ _01351_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__o21a_1
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6559_ MuI._2449_ MuI._2455_ MuI._2442_ MuI._2446_ vssd1 vssd1 vccd1 vccd1 MuI._2458_
+ sky130_fd_sc_hd__o211a_1
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5778__A MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__A1 _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _02096_ _02194_ _05176_ net17 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__and4_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07868__B2 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _00077_ _04369_ vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__nand2_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08596_ _01203_ _01211_ _01213_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__and3_1
XFILLER_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__A2 _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _00162_ _05638_ _00163_ _00164_ vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12613__A1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07478_ net117 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _01831_ _01796_ _01833_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__or4_2
XANTENNA__11611__B _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__C _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13169__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07089__A _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__A2 _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _01762_ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and2b_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11330__C _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6121__B MuI._1975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10227__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _06545_ _00059_ _01682_ _01681_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a31o_1
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3518__A1 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _03860_ _03738_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__or2_2
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12090_ _04777_ _04782_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__and2_1
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06721__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12442__B _05198_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3761__A MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _00414_ _06622_ net130 net129 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__and4_1
XANTENNA__08348__A2 _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._533__B1 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _03615_ _05660_ _05883_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21boi_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10897__B _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input13_A a_operand[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13273__B _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ _04757_ _04758_ _04604_ _04610_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__o211a_1
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _00095_ net117 _06466_ _06461_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__and4_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _03551_ _03552_ _03368_ _03535_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__a211oi_1
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ _03280_ _03283_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__nand2_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11521__B _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ _06387_ _06389_ _04635_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__mux2_1
X_10687_ _03205_ _03203_ _03204_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10418__A _03113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3757__A1 MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12426_ _00088_ _03247_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nand2_1
XFILLER_173_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5930_ MuI._1460_ MuI._1645_ MuI._1761_ MuI._1763_ MuI._1765_ vssd1 vssd1 vccd1
+ vccd1 MuI._1766_ sky130_fd_sc_hd__o311a_1
XFILLER_154_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11040__B1 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12357_ _00506_ _00676_ _06525_ _06568_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__and4_1
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._810_ AuI.pe.significand\[14\] AuI.pe.significand\[15\] AuI.pe._367_ AuI.pe.significand\[13\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._349_ sky130_fd_sc_hd__or4b_1
XANTENNA__07795__B1 _05380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5861_ MuI._1614_ MuI._1616_ MuI._1617_ vssd1 vssd1 vccd1 vccd1 MuI._1690_ sky130_fd_sc_hd__o21ba_1
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output81_A net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _00462_ _06518_ _06562_ _00086_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07727__A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _05128_ _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nand2_1
XFILLER_206_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4812_ MuI._0532_ MuI._0534_ MuI._0535_ vssd1 vssd1 vccd1 vccd1 MuI._0536_ sky130_fd_sc_hd__a21oi_1
XAuI.pe._741_ AuI.pe._380_ AuI.pe._389_ AuI.pe._390_ vssd1 vssd1 vccd1 vccd1 AuI.pe._286_
+ sky130_fd_sc_hd__a21o_1
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5792_ MuI._2451_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._1614_ sky130_fd_sc_hd__nand2_1
XANTENNA__09536__B2 _02078_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10153__A _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1666_ AuI._0018_ vssd1 vssd1 vccd1 vccd1 AuI.result\[28\] sky130_fd_sc_hd__clkbuf_1
X_11239_ _03859_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._672_ AuI.pe._145_ AuI.pe._002_ AuI.pe._053_ AuI.pe._158_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._221_ sky130_fd_sc_hd__a22o_1
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07547__B1 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4743_ MuI._0457_ MuI._0459_ vssd1 vssd1 vccd1 vccd1 MuI._0461_ sky130_fd_sc_hd__or2_1
XANTENNA__12540__B1 _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._1597_ AuI.pe.Significand\[13\] AuI._0769_ vssd1 vssd1 vccd1 vccd1 AuI._0770_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4674_ MuI._0380_ MuI._0384_ vssd1 vssd1 vccd1 vccd1 MuI._0385_ sky130_fd_sc_hd__and2b_1
XFILLER_95_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ _03056_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__buf_6
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6413_ MuI._2151_ MuI._2152_ vssd1 vssd1 vccd1 vccd1 MuI._2298_ sky130_fd_sc_hd__and2_1
XMuI._3625_ MuI._2176_ MuI._2187_ vssd1 vssd1 vccd1 vccd1 MuI._2231_ sky130_fd_sc_hd__xor2_1
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07462__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6344_ MuI._3091_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._2222_ sky130_fd_sc_hd__nand2_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3556_ MuI._1461_ vssd1 vssd1 vccd1 vccd1 MuI._1472_ sky130_fd_sc_hd__buf_2
XFILLER_35_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08450_ _02840_ _04531_ _01031_ _01030_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._5434__A1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__C _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5434__B2 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5748__D MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._827__A1 AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6275_ MuI._2074_ MuI._2101_ MuI._2073_ vssd1 vssd1 vccd1 vccd1 MuI._2146_ sky130_fd_sc_hd__a21boi_1
X_07401_ _00016_ _00017_ _00018_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__a21o_1
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3487_ MuI._0691_ MuI._0548_ MuI._0702_ vssd1 vssd1 vccd1 vccd1 MuI._0713_ sky130_fd_sc_hd__o21a_1
XANTENNA__13399__A2 _06305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08381_ _00996_ _00997_ _00998_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__and3_1
XFILLER_177_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12808__A _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5226_ MuI._0990_ MuI._0991_ vssd1 vssd1 vccd1 vccd1 MuI._0992_ sky130_fd_sc_hd__nor2_1
XFILLER_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07332_ _06598_ _06599_ _04896_ _04961_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__and4_1
XFILLER_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06806__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5157_ MuI._2429_ MuI._3402_ MuI._3396_ MuI._2660_ vssd1 vssd1 vccd1 vccd1 MuI._0916_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11431__B _04076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ net107 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__buf_4
XFILLER_177_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0874__A1 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4108_ MuI._2798_ MuI._3207_ vssd1 vssd1 vccd1 vccd1 MuI._3208_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _01415_ _01435_ _01434_ _01431_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__o211ai_1
XMuI._5088_ MuI._0838_ MuI._0839_ vssd1 vssd1 vccd1 vccd1 MuI._0840_ sky130_fd_sc_hd__or2b_1
XFILLER_192_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07194_ net116 vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__buf_4
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4039_ MuI._3135_ MuI._3138_ vssd1 vssd1 vccd1 vccd1 MuI._3139_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12543__A _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6162__A2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _02544_ _02554_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__nor3_1
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__A _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10063__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A a_operand[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _02404_ _02405_ _02487_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11309__D _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5633__A1_N MuI._3269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09766_ _02361_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__nand3_1
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06978_ _05187_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08468__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08717_ _01333_ _01334_ _06475_ _00040_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__and4bb_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12834__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _02088_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__xor2_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__B2 _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _01168_ _01265_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__or2_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6116__B MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _01195_ _01194_ _01187_ _01193_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__o211ai_2
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__A _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ _04068_ _02259_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2b_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _04376_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06716__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10073__A1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3756__A MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ _06560_ _05649_ _03246_ _03248_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a22o_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ _02827_ _02875_ _06108_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__o21ai_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ _03172_ _03173_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__nor2_1
XFILLER_182_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12211_ _04909_ _04911_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nor2_1
XFILLER_151_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ _06095_ _06096_ _02925_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__mux2_1
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__A2 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _04839_ _04844_ _04970_ _04971_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a211oi_2
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3491__A MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1520_ AuI._0704_ AuI._0654_ vssd1 vssd1 vccd1 vccd1 AuI._0705_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07266__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12073_ _02844_ _04892_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__o21a_1
XFILLER_110_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09184__D _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ _03764_ _03765_ _03767_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21o_1
XAuI._1451_ AuI._0422_ AuI._0439_ AuI._0444_ vssd1 vssd1 vccd1 vccd1 AuI._0637_ sky130_fd_sc_hd__a21o_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1382_ AuI._0569_ AuI._0573_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[20\]
+ sky130_fd_sc_hd__xnor2_4
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4467__A2 MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10701__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07282__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11089__B1 _02711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12286__C1 _05127_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12975_ _05603_ _05782_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__nor2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6307__A MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10420__B _00811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4390_ MuI._0071_ MuI._0072_ vssd1 vssd1 vccd1 vccd1 MuI._0073_ sky130_fd_sc_hd__and2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _04738_ _04739_ _04722_ _04587_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__o211ai_1
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _00221_ _05660_ _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a22o_1
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12628__A _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6060_ MuI._3154_ MuI._1842_ MuI._1908_ vssd1 vssd1 vccd1 vccd1 MuI._1909_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _03165_ _03169_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a211oi_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09454__B1 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5011_ MuI._0751_ MuI._0752_ vssd1 vssd1 vccd1 vccd1 MuI._0755_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ _04589_ _04590_ _04570_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__a21o_1
XFILLER_159_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3666__A MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10739_ _03254_ _03255_ _03264_ _03263_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a31o_1
XFILLER_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _06304_ _02699_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nor2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08841__A _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09477__A1_N _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._588__A3 AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _02752_ _05142_ _05143_ _05259_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__a31o_4
XANTENNA__11013__B1 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ _02817_ _05883_ _06258_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__nand3b_1
XANTENNA__12363__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__B1 _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5913_ MuI._1743_ MuI._1744_ MuI._1745_ vssd1 vssd1 vccd1 vccd1 MuI._1748_ sky130_fd_sc_hd__nand3_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5844_ MuI.b_operand\[11\] MuI._0088_ MuI._0694_ MuI._0695_ vssd1 vssd1 vccd1
+ vccd1 MuI._1672_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13305__A2 _06208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _03002_ _04520_ _00045_ _00050_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__o2bb2a_1
XAuI.pe._724_ AuI.pe._211_ AuI.pe._208_ AuI.pe.significand\[20\] AuI.pe._076_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._270_ sky130_fd_sc_hd__or4b_1
XMuI._5775_ MuI._1591_ MuI._1592_ MuI._1594_ vssd1 vssd1 vccd1 vccd1 MuI._1596_ sky130_fd_sc_hd__a21oi_1
X_06901_ _04358_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._5105__B MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1649_ AuI.exponent_sub\[2\] AuI._0695_ AuI._0602_ AuI._0719_ AuI._0699_ vssd1
+ vssd1 vccd1 vccd1 AuI._0005_ sky130_fd_sc_hd__o221a_1
X_07881_ _00497_ _00498_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__or2_1
XFILLER_68_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._655_ AuI.pe._105_ AuI.pe._086_ AuI.pe._200_ AuI.pe._204_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._205_ sky130_fd_sc_hd__a211o_1
XFILLER_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4726_ MuI._0878_ MuI._0112_ MuI._0308_ vssd1 vssd1 vccd1 vccd1 MuI._0442_ sky130_fd_sc_hd__a21oi_1
X_09620_ _02204_ _02207_ _02206_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a21o_1
XANTENNA__11707__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06832_ _03615_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4657_ MuI._0253_ MuI._0365_ vssd1 vssd1 vccd1 vccd1 MuI._0366_ sky130_fd_sc_hd__or2_1
XAuI.pe._586_ AuI.pe._140_ vssd1 vssd1 vccd1 vccd1 AuI.pe._141_ sky130_fd_sc_hd__clkbuf_2
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09551_ _02177_ _02181_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a21oi_1
XFILLER_83_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06763_ _02873_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[14\] sky130_fd_sc_hd__clkbuf_4
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10330__B _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3608_ MuI._2022_ MuI._2033_ vssd1 vssd1 vccd1 vccd1 MuI._2044_ sky130_fd_sc_hd__or2_1
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08502_ _01007_ _01051_ _01052_ _01053_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__a211o_1
XFILLER_64_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4588_ MuI._2473_ MuI._2830_ MuI._0216_ MuI._0217_ vssd1 vssd1 vccd1 vccd1 MuI._0290_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06694_ _02129_ net1 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__and2_1
X_09482_ _02091_ _02093_ _02092_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10171__A_N _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07342__D net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3539_ MuI._1274_ vssd1 vssd1 vccd1 vccd1 MuI._1285_ sky130_fd_sc_hd__clkbuf_4
XMuI._6327_ MuI._2178_ vssd1 vssd1 vccd1 vccd1 MuI._2203_ sky130_fd_sc_hd__inv_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08433_ _01007_ _01008_ _01014_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__nand3_1
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6258_ MuI._0790_ MuI._1274_ vssd1 vssd1 vccd1 vccd1 MuI._2127_ sky130_fd_sc_hd__nand2_1
XFILLER_51_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08364_ _00978_ _00981_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5209_ MuI._0883_ MuI._0884_ MuI._0894_ vssd1 vssd1 vccd1 vccd1 MuI._0973_ sky130_fd_sc_hd__and3_1
XANTENNA__12257__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6189_ MuI._2939_ MuI._2811_ MuI._2843_ MuI._2840_ vssd1 vssd1 vccd1 vccd1 MuI._2051_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11252__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _06597_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and2_1
XANTENNA__08799__A2 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ _00728_ _00727_ _04046_ _00303_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__and4_1
XANTENNA__09269__D net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__D net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ _06545_ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nand2_1
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ _06475_ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__nand2_1
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A2 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5894__A1 MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._494__A AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__B1 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5894__B2 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12720__B _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09818_ _02442_ _03884_ _02455_ _02456_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__a211oi_1
XFILLER_98_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11617__A _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09749_ _02342_ _02323_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__and2_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07533__C net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ _05513_ _05516_ _05514_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__o21ba_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11711_ _04505_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__xnor2_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12691_ _05559_ _05560_ _05435_ _05491_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__a211o_1
XFILLER_187_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _02965_ _04725_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__nand2_1
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _04302_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__inv_2
XFILLER_211_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 a_operand[21] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_6
X_13312_ _02830_ _06220_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__nand2_1
X_10524_ _03227_ _03229_ _03230_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a21o_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 a_operand[31] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_8
XFILLER_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0951_ AuI._0154_ AuI._0162_ vssd1 vssd1 vccd1 vccd1 AuI._0163_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _02837_ _06150_ _06082_ _02711_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a31o_1
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0882_ AuI._0096_ AuI._0097_ AuI._0100_ AuI._0101_ vssd1 vssd1 vccd1 vccd1 AuI._0102_
+ sky130_fd_sc_hd__or4_1
X_10455_ _03798_ _04133_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__nand2_1
XFILLER_183_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11546__B2 _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07277__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13174_ _02841_ _06075_ _06077_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__nand4_1
X_10386_ _00164_ _00162_ _00783_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand4_1
XFILLER_112_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__A_N _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3890_ MuI._2911_ MuI._2912_ vssd1 vssd1 vccd1 vccd1 MuI._2990_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._4748__C MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12125_ _04951_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__xor2_2
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13299__B2 _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07427__D _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1503_ AuI._0583_ AuI._0586_ vssd1 vssd1 vccd1 vccd1 AuI._0689_ sky130_fd_sc_hd__nor2_1
X_12056_ _02575_ _02579_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and2_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6736__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12630__B _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5560_ MuI._1344_ MuI._1345_ MuI._1357_ vssd1 vssd1 vccd1 vccd1 MuI._1359_ sky130_fd_sc_hd__and3_1
X_11007_ _03562_ _03564_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1434_ AuI._0617_ AuI._0619_ vssd1 vssd1 vccd1 vccd1 AuI._0620_ sky130_fd_sc_hd__or2_1
XFILLER_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4511_ MuI._0181_ MuI._0182_ vssd1 vssd1 vccd1 vccd1 MuI._0205_ sky130_fd_sc_hd__nor2_1
XAuI.pe._440_ AuI.pe._399_ AuI.pe._002_ AuI.pe._004_ AuI.pe._006_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._007_ sky130_fd_sc_hd__or4_1
XFILLER_93_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10521__A2 _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5491_ MuI._1227_ MuI._1281_ MuI._1272_ MuI._1280_ vssd1 vssd1 vccd1 vccd1 MuI._1283_
+ sky130_fd_sc_hd__a211o_1
XAuI._1365_ AuI._0539_ AuI._0540_ AuI._0546_ AuI._0557_ vssd1 vssd1 vccd1 vccd1 AuI._0558_
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07443__C _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10150__B _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4442_ MuI._3390_ MuI._3421_ vssd1 vssd1 vccd1 vccd1 MuI._0129_ sky130_fd_sc_hd__xor2_1
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _05338_ _02745_ _02722_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a21o_1
XAuI._1296_ AuI._0257_ AuI._0491_ AuI._0492_ AuI._0493_ vssd1 vssd1 vccd1 vccd1 AuI._0495_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4373_ MuI._2660_ MuI._2440_ MuI._2844_ MuI._2845_ vssd1 vssd1 vccd1 vccd1 MuI._0055_
+ sky130_fd_sc_hd__and4_1
XFILLER_179_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ _04572_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nand3_1
XFILLER_178_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6112_ MuI._2851_ MuI._0526_ MuI._1887_ MuI._1965_ vssd1 vssd1 vccd1 vccd1 MuI._1966_
+ sky130_fd_sc_hd__a31oi_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _02809_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__or2_1
XANTENNA__07150__A1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6043_ MuI._1886_ MuI._1889_ vssd1 vssd1 vccd1 vccd1 MuI._1891_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3820__B1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07100_ _06413_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _00693_ _00696_ _00697_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__nand3_2
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07031_ _05756_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__clkbuf_4
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12093__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__A1 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07187__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6876_ MuI._2775_ MuI._2500_ vssd1 vssd1 vccd1 vccd1 MuI._2776_ sky130_fd_sc_hd__xnor2_1
XFILLER_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08982_ _01335_ _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__nor2_1
XMuI._5827_ MuI._1285_ MuI._0321_ MuI._1562_ MuI._1561_ vssd1 vssd1 vccd1 vccd1 MuI._1653_
+ sky130_fd_sc_hd__a31o_1
X_07933_ _06620_ _00550_ _06582_ _06586_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_AuI._1006__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4955__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._707_ AuI.pe._244_ AuI.pe._245_ AuI.pe._252_ AuI.pe._253_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._254_ sky130_fd_sc_hd__or4_1
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08166__B1 _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5758_ MuI._2854_ MuI._2341_ MuI._0085_ MuI._2853_ vssd1 vssd1 vccd1 vccd1 MuI._1577_
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07864_ _00360_ _00365_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__or2b_1
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._638_ AuI.pe._393_ AuI.pe._399_ AuI.pe._002_ AuI.pe._380_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._189_ sky130_fd_sc_hd__a22o_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07913__B1 _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4709_ MuI._2693_ MuI._2638_ MuI._3349_ MuI._0088_ vssd1 vssd1 vccd1 vccd1 MuI._0423_
+ sky130_fd_sc_hd__and4_1
X_09603_ _02202_ _02201_ _02193_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a21o_1
XFILLER_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06815_ _03432_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__buf_4
XMuI._5689_ MuI._1498_ MuI._1499_ MuI._1482_ vssd1 vssd1 vccd1 vccd1 MuI._1501_ sky130_fd_sc_hd__a21o_1
X_07795_ _06682_ _00412_ _05380_ _00000_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a22oi_2
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._569_ AuI.pe._380_ vssd1 vssd1 vccd1 vccd1 AuI.pe._125_ sky130_fd_sc_hd__clkbuf_4
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _02161_ _02163_ _02090_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08168__D _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06746_ _02691_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[10\] sky130_fd_sc_hd__buf_2
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13462__A1 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07650__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _02069_ _02074_ _02087_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__or3_1
XFILLER_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11172__A _00414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08416_ _01027_ _01028_ _01033_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__nand3_2
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._120_ FuI._050_ FuI._056_ FuI._024_ FuI._030_ FuI.a_operand\[16\] vssd1 vssd1
+ vccd1 vccd1 FuI._006_ sky130_fd_sc_hd__o311a_1
X_09396_ _02003_ _02008_ _02012_ _02013_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__o211ai_2
XFILLER_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4603__A2 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08347_ _06475_ _00534_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__nand2_1
XFILLER_193_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _00894_ _00895_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__or2_2
XANTENNA__08481__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07229_ _06526_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07097__A _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10240_ _02775_ _02811_ _02874_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o31a_2
XFILLER_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__B _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _03024_ _05058_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__and2b_1
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10950__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08157__B1 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10889__C _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4584__B MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._488__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ _05690_ _05691_ _00077_ _05831_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__and4bb_1
XAuI._1150_ AuI._0212_ AuI._0351_ AuI._0354_ AuI._0357_ AuI._0249_ vssd1 vssd1 vccd1
+ vccd1 AuI._0358_ sky130_fd_sc_hd__a311o_2
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09657__B1 _00072_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12256__A2 _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10267__A1 _00672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _00283_ _03071_ _05616_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a22o_1
XAuI._1081_ AuI._0199_ AuI._0200_ AuI._0201_ vssd1 vssd1 vccd1 vccd1 AuI._0292_ sky130_fd_sc_hd__and3_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08375__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11082__A _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12674_ _05455_ _05458_ _05543_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__o211ai_2
XANTENNA__08806__D _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4750__D MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ _04405_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__xor2_1
XFILLER_168_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11556_ _03134_ _04323_ _04324_ _04336_ _04342_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__a311o_2
XANTENNA__12625__B _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _03202_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0934_ AuI._0130_ AuI._0131_ AuI._0144_ AuI._0145_ vssd1 vssd1 vccd1 vccd1 AuI._0146_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07719__B _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10426__A _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ _00502_ _04542_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4759__B MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ _06029_ _06032_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__a21o_1
XMuI._4991_ MuI._0725_ MuI._0726_ MuI._0732_ vssd1 vssd1 vccd1 vccd1 MuI._0733_ sky130_fd_sc_hd__or3_1
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ _02999_ _02998_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__or2b_1
XFILLER_124_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0865_ AuI._0079_ AuI._0081_ AuI._0083_ AuI._0084_ vssd1 vssd1 vccd1 vccd1 AuI._0085_
+ sky130_fd_sc_hd__or4_1
XANTENNA__10145__B _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6730_ MuI._2645_ vssd1 vssd1 vccd1 vccd1 MuI._2646_ sky130_fd_sc_hd__clkinv_2
XFILLER_124_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3942_ MuI._0768_ MuI._2836_ MuI._2845_ MuI._0559_ vssd1 vssd1 vccd1 vccd1 MuI._3042_
+ sky130_fd_sc_hd__a22oi_2
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _06058_ _06060_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__and2_1
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10369_ _03061_ _03062_ _03044_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21oi_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3873_ MuI._1472_ MuI._2841_ vssd1 vssd1 vccd1 vccd1 MuI._2973_ sky130_fd_sc_hd__nand2_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6661_ MuI._1837_ MuI._2569_ vssd1 vssd1 vccd1 vccd1 MuI._2570_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12108_ _04803_ _04785_ _04784_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a21boi_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _05986_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__or2_1
XMuI._5612_ MuI._3397_ MuI._0112_ MuI._0246_ MuI._3403_ vssd1 vssd1 vccd1 vccd1 MuI._1416_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6592_ MuI._0262_ MuI._0251_ MuI._0229_ vssd1 vssd1 vccd1 vccd1 MuI._2494_ sky130_fd_sc_hd__and3b_1
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12039_ _04766_ _04746_ _04860_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a211o_2
XFILLER_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4494__B MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5543_ MuI._1335_ MuI._1339_ MuI._2876_ MuI._0321_ vssd1 vssd1 vccd1 vccd1 MuI._1341_
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1417_ AuI.operand_a\[26\] AuI.operand_a\[27\] AuI._0603_ vssd1 vssd1 vccd1 vccd1
+ AuI._0604_ sky130_fd_sc_hd__and3_1
XFILLER_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._423_ AuI.pe.significand\[15\] AuI.pe.significand\[14\] vssd1 vssd1 vccd1
+ vccd1 AuI.pe._390_ sky130_fd_sc_hd__and2b_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._5474_ MuI._1261_ MuI._1264_ vssd1 vssd1 vccd1 vccd1 MuI._1265_ sky130_fd_sc_hd__xor2_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5102__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1348_ AuI._0538_ AuI._0541_ AuI._0542_ vssd1 vssd1 vccd1 vccd1 AuI._0543_ sky130_fd_sc_hd__and3_1
X_07580_ _06610_ _00197_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__nand2_1
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4425_ MuI._0110_ vssd1 vssd1 vccd1 vccd1 MuI._0111_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07470__A net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11704__B _00878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1279_ AuI._0455_ AuI._0456_ AuI._0468_ AuI._0469_ vssd1 vssd1 vccd1 vccd1 AuI._0479_
+ sky130_fd_sc_hd__and4_1
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08320__B1 _00617_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4356_ MuI._3395_ MuI._3406_ vssd1 vssd1 vccd1 vccd1 MuI._0036_ sky130_fd_sc_hd__xnor2_2
XFILLER_179_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _01659_ _01661_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nand2_1
XFILLER_33_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ _00632_ _00629_ _00631_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__nand3_1
XMuI._4287_ MuI._3382_ MuI._3386_ vssd1 vssd1 vccd1 vccd1 MuI._3387_ sky130_fd_sc_hd__nand2_1
XFILLER_194_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _01784_ _01796_ _01797_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__nor3_1
XFILLER_175_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6026_ MuI._1870_ MuI._1871_ vssd1 vssd1 vccd1 vccd1 MuI._1872_ sky130_fd_sc_hd__nor2_1
XFILLER_159_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12955__B1 _04211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08132_ _00394_ _00403_ _00402_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a21o_1
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06814__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3854__A MuI._2926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08063_ _06439_ _00303_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__nand2_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6230__A MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout113_A net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09547__D _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07014_ _05574_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_134_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12183__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6859_ MuI._2490_ MuI._2488_ vssd1 vssd1 vccd1 vccd1 MuI._2762_ sky130_fd_sc_hd__or2b_1
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08965_ _01578_ _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11167__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _06623_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__clkbuf_8
XFILLER_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08896_ _06578_ _02647_ _04574_ _00030_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__and4_1
XANTENNA__12486__A2 _04994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ _00461_ _00463_ _00464_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__or3_1
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13435__A1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07778_ _06663_ _06666_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__nand2_1
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08476__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07380__A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09517_ _01981_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__and3_1
X_06729_ _02507_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08195__B _00812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4037__B1 MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ _02069_ _02070_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__or2_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._103_ net104 FuI.a_operand\[23\] vssd1 vssd1 vccd1 vccd1 FuI._061_ sky130_fd_sc_hd__and2_1
X_09379_ net68 net38 net126 net125 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__and4_1
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08923__B _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ _04052_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__inv_2
X_12390_ _05126_ _05128_ _05236_ _05237_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__a211oi_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__A _01714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _04107_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__xor2_4
XFILLER_181_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11272_ _06585_ _06583_ _00785_ _00153_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__and4_1
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4760__A1 MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _05782_ _05903_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__or2_1
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10223_ _02807_ _02906_ _02806_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4760__B2 MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12461__A _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input43_A b_operand[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _03507_ _05671_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ _04251_ _02388_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__and2b_1
XFILLER_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09770__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11685__B1 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1202_ AuI._0276_ AuI._0405_ AuI._0406_ vssd1 vssd1 vccd1 vccd1 AuI._0407_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11805__A _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__A _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1133_ AuI._0334_ AuI._0249_ AuI._0341_ vssd1 vssd1 vccd1 vccd1 AuI._0342_ sky130_fd_sc_hd__or3b_2
XFILLER_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4210_ MuI._3308_ MuI._3309_ vssd1 vssd1 vccd1 vccd1 MuI._3310_ sky130_fd_sc_hd__or2_1
X_10987_ _03725_ _03726_ _03715_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5190_ MuI._0928_ MuI._0929_ MuI._0950_ MuI._0951_ vssd1 vssd1 vccd1 vccd1 MuI._0952_
+ sky130_fd_sc_hd__and4bb_1
XANTENNA_MuI._4761__C MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _05525_ _05526_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or2_1
XAuI._1064_ AuI._0265_ AuI._0268_ AuI._0271_ AuI._0273_ AuI._0274_ AuI._0209_ vssd1
+ vssd1 vccd1 vccd1 AuI._0275_ sky130_fd_sc_hd__mux4_1
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4141_ MuI._3236_ MuI._3240_ vssd1 vssd1 vccd1 vccd1 MuI._3241_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4480__D MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ net61 _05209_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__nand2_1
XFILLER_157_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12636__A _00299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__B _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4072_ MuI._3160_ MuI._3171_ vssd1 vssd1 vccd1 vccd1 MuI._3172_ sky130_fd_sc_hd__nand2_1
XFILLER_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _04395_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nand3_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12401__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12588_ _05449_ _05450_ _05446_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__a21o_1
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ _04322_ _04312_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__or2b_1
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10156__A _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0917_ net23 net55 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0134_ sky130_fd_sc_hd__mux2_1
XFILLER_125_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13467__A _06376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ _03755_ _05713_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__nand3_1
XMuI._4974_ MuI._1263_ MuI._0445_ MuI._0622_ MuI._0623_ vssd1 vssd1 vccd1 vccd1 MuI._0715_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._0848_ net121 vssd1 vssd1 vccd1 vccd1 AuI._0068_ sky130_fd_sc_hd__inv_2
XFILLER_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6713_ MuI._2387_ MuI._2623_ MuI._2337_ vssd1 vssd1 vccd1 vccd1 MuI._2628_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11912__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3925_ MuI._3020_ MuI._3024_ vssd1 vssd1 vccd1 vccd1 MuI._3025_ sky130_fd_sc_hd__xor2_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07465__A _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6644_ MuI._1458_ MuI._1238_ vssd1 vssd1 vccd1 vccd1 MuI._2552_ sky130_fd_sc_hd__and2b_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3856_ MuI._2944_ MuI._2943_ vssd1 vssd1 vccd1 vccd1 MuI._2956_ sky130_fd_sc_hd__and2b_1
X_08750_ _01366_ _01367_ _06680_ _00074_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__and4bb_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07701_ _00288_ _00293_ vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__or2_1
XFILLER_78_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3787_ MuI._0482_ MuI._0493_ MuI._2886_ vssd1 vssd1 vccd1 vccd1 MuI._2887_ sky130_fd_sc_hd__a21bo_1
XMuI._6575_ MuI._1648_ MuI._1714_ MuI._1736_ vssd1 vssd1 vccd1 vccd1 MuI._2476_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._5113__B MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08681_ _01297_ _01296_ _01295_ _01291_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__o211a_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07344__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5526_ MuI._1260_ MuI._1268_ MuI._1267_ vssd1 vssd1 vccd1 vccd1 MuI._1322_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07344__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__B1 _04176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _00247_ _00248_ _00020_ _00021_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__o211ai_1
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._406_ AuI.pe.significand\[9\] AuI.pe.significand\[10\] AuI.pe.significand\[11\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._373_ sky130_fd_sc_hd__or3_1
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06809__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5457_ MuI._3306_ MuI._3307_ MuI.a_operand\[4\] MuI.a_operand\[3\] vssd1 vssd1
+ vccd1 vccd1 MuI._1246_ sky130_fd_sc_hd__and4_1
XFILLER_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07563_ _00178_ _00179_ _00174_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__a21o_1
XANTENNA__11434__B _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4408_ MuI._0087_ MuI._0090_ MuI._0091_ vssd1 vssd1 vccd1 vccd1 MuI._0092_ sky130_fd_sc_hd__o21ai_1
X_09302_ _01805_ _01801_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5388_ MuI._1160_ MuI._1168_ MuI._1169_ vssd1 vssd1 vccd1 vccd1 MuI._1170_ sky130_fd_sc_hd__or3b_1
XFILLER_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07494_ _00109_ _00110_ _00111_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__or3_1
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4339_ MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 MuI._0017_ sky130_fd_sc_hd__buf_2
XFILLER_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09233_ _01644_ _01645_ _01661_ _01662_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and4bb_1
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09839__B _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12546__A _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ _01780_ _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or2b_1
XMuI._6009_ MuI._1274_ MuI._2849_ vssd1 vssd1 vccd1 vccd1 MuI._1853_ sky130_fd_sc_hd__nand2_1
XFILLER_175_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08115_ _00731_ _00732_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10066__A _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ _01368_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4399__B MuI._2374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08046_ _00662_ _00661_ _00528_ _00527_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__o211ai_4
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4742__A1 MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__B1 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10706__A2 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10105__A_N _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09997_ _01316_ _01275_ _01315_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__and3_1
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5298__A2 MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13105__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08780__B1 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4846__C MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08948_ _01508_ _01532_ _01564_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__o211a_1
XFILLER_57_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08879_ _02539_ _04660_ _01476_ _01475_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__a31o_1
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__A2 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08532__B1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _03643_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__xnor2_2
XFILLER_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _04698_ _04699_ _04662_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4862__B MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08637__C _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ _03568_ _03569_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nand3_4
XANTENNA__10890__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10890__B2 _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08884__A2_N _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__B1 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10772_ MuI.result\[3\] _02737_ _06045_ FuI.Integer\[3\] vssd1 vssd1 vccd1 vccd1
+ _03498_ sky130_fd_sc_hd__a22o_1
XFILLER_201_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12511_ _02621_ _05368_ _02619_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a21oi_2
XFILLER_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5758__B1 MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ _06404_ _06405_ _06363_ _06406_ _03134_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__o311a_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5222__A2 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _06439_ _05198_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__nand2_1
XANTENNA__09468__C net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08899__A2_N _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3494__A MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _05182_ _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nor3_4
XFILLER_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ _04052_ _04053_ _04090_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o22a_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4102__B MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13344__B1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ AuI.result\[6\] _02731_ _04018_ _02935_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__a22o_1
XFILLER_107_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10704__A _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _02496_ _04391_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and2b_1
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3941__B MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11186_ _03941_ _03942_ _03919_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3710_ MuI._2783_ MuI._2784_ MuI._2808_ vssd1 vssd1 vccd1 vccd1 MuI._2810_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4690_ MuI._0183_ MuI._0204_ vssd1 vssd1 vccd1 vccd1 MuI._0402_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09123__A1_N _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08771__B1 _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _02812_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__and2b_1
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3641_ MuI.b_operand\[22\] MuI.b_operand\[21\] MuI._2363_ vssd1 vssd1 vccd1 vccd1
+ MuI._2407_ sky130_fd_sc_hd__and3_1
XFILLER_208_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__buf_6
XANTENNA_MuI._6238__A1 MuI._0350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6238__B2 MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6360_ MuI._2194_ MuI._2199_ MuI._2237_ MuI._2238_ vssd1 vssd1 vccd1 vccd1 MuI._2239_
+ sky130_fd_sc_hd__a211oi_1
XMuI._3572_ MuI._1593_ MuI._1615_ MuI._1637_ vssd1 vssd1 vccd1 vccd1 MuI._1648_ sky130_fd_sc_hd__nand3_1
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5311_ MuI._0964_ MuI._0961_ MuI._0963_ vssd1 vssd1 vccd1 vccd1 MuI._1085_ sky130_fd_sc_hd__nand3_1
XFILLER_211_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6291_ MuI._2127_ MuI._2129_ MuI._2128_ vssd1 vssd1 vccd1 vccd1 MuI._2163_ sky130_fd_sc_hd__o21ba_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09079__A1 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5242_ MuI._0993_ MuI._0994_ MuI._1008_ vssd1 vssd1 vccd1 vccd1 MuI._1009_ sky130_fd_sc_hd__a21o_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1116_ AuI._0324_ AuI._0325_ vssd1 vssd1 vccd1 vccd1 AuI._0326_ sky130_fd_sc_hd__and2_2
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08844__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5173_ MuI._2853_ MuI._2854_ MuI._0100_ MuI._3245_ vssd1 vssd1 vccd1 vccd1 MuI._0934_
+ sky130_fd_sc_hd__and4_1
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _02856_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or2b_1
XFILLER_176_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1047_ AuI._0258_ vssd1 vssd1 vccd1 vccd1 AuI._0259_ sky130_fd_sc_hd__buf_2
XMuI._4124_ MuI._3000_ MuI._2754_ MuI._2790_ MuI._3223_ vssd1 vssd1 vccd1 vccd1 MuI._3224_
+ sky130_fd_sc_hd__and4_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4421__B1 MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4055_ MuI._3153_ MuI._3081_ MuI._3084_ vssd1 vssd1 vccd1 vccd1 MuI._3155_ sky130_fd_sc_hd__and3_1
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08054__A2 _00518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._587__A AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07262__B1 _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _02444_ _02446_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__and2_1
XFILLER_160_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07195__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4957_ MuI._0694_ MuI._0695_ MuI.b_operand\[11\] MuI._0088_ vssd1 vssd1 vccd1
+ vccd1 MuI._0696_ sky130_fd_sc_hd__and4bb_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09851_ _02500_ _02497_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__xnor2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11429__B _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3908_ MuI._3006_ MuI._3007_ vssd1 vssd1 vccd1 vccd1 MuI._3008_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._4666__C MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08802_ _00444_ _06437_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nand2_2
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4888_ MuI._2473_ MuI._3372_ MuI._0430_ MuI._0431_ vssd1 vssd1 vccd1 vccd1 MuI._0620_
+ sky130_fd_sc_hd__o2bb2a_1
X_09782_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__nor2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ net19 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6627_ MuI._2527_ MuI._2529_ MuI._2532_ vssd1 vssd1 vccd1 vccd1 MuI._2533_ sky130_fd_sc_hd__a21o_1
XFILLER_100_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3839_ MuI.b_operand\[19\] vssd1 vssd1 vccd1 vccd1 MuI._2939_ sky130_fd_sc_hd__buf_2
X_08733_ _02647_ _00084_ _04574_ _02582_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__a22o_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._542__B2 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__C _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6558_ MuI._2456_ vssd1 vssd1 vccd1 vccd1 MuI._2457_ sky130_fd_sc_hd__inv_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08664_ _06495_ _05176_ _05241_ _02107_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__a22oi_2
XFILLER_82_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5778__B MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07868__A2 _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5509_ MuI._1255_ MuI._1253_ MuI._1254_ vssd1 vssd1 vccd1 vccd1 MuI._1303_ sky130_fd_sc_hd__or3_1
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07615_ _00093_ _00230_ _00232_ vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__a21bo_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6489_ MuI._2375_ MuI._2372_ vssd1 vssd1 vccd1 vccd1 MuI._2381_ sky130_fd_sc_hd__xor2_2
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _01171_ _01212_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__and2b_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07546_ _06479_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__buf_4
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5794__A MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11821__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07477_ net118 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__buf_2
XFILLER_195_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09216_ _01830_ _01829_ _01828_ _01825_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__o211a_1
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08904__D _00083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__C _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09147_ _01762_ _01763_ _01764_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__or3_1
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._497__A AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09078_ _01680_ _01694_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nand3_2
XANTENNA_MuI._3518__A2 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08029_ _06641_ _00645_ _00644_ _00641_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__a211o_1
XFILLER_123_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ _06583_ _06537_ _05756_ _06585_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a22oi_2
XANTENNA_AuI.pe._781__A1 AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4479__B1 MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12991_ _03550_ _03449_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nand2_2
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _04755_ _04756_ _04652_ _04653_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o211a_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _00462_ _05498_ _05563_ _00237_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__a22oi_2
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _03368_ _03535_ _03551_ _03552_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__o211a_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10755_ _03334_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__xnor2_2
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ _06364_ _06388_ _02918_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a21o_1
XANTENNA__11521__C _04303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ _03403_ _03401_ _03402_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand3_1
XFILLER_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10418__B _03116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3757__A2 MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ _00237_ _00462_ _00785_ _00153_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__and4_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11040__A1 _06583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11040__B2 _06585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _06442_ _00002_ _06561_ _06444_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__a22oi_1
XANTENNA__06912__A _04467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07795__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5860_ MuI._1599_ MuI._1601_ MuI._1600_ vssd1 vssd1 vccd1 vccd1 MuI._1689_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__A _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _05126_ _05127_ _05033_ _05034_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a211o_1
XAuI.pe._740_ AuI.pe._211_ AuI.pe._000_ AuI.pe._384_ AuI.pe._042_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._285_ sky130_fd_sc_hd__a31o_1
XFILLER_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4811_ MuI._0529_ MuI._0531_ vssd1 vssd1 vccd1 vccd1 MuI._0535_ sky130_fd_sc_hd__and2b_1
XANTENNA_output74_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5791_ MuI._1609_ MuI._1611_ MuI._1610_ vssd1 vssd1 vccd1 vccd1 MuI._1613_ sky130_fd_sc_hd__a21o_1
X_11238_ _03997_ _03999_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__xnor2_4
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1665_ AuI._0015_ AuI._0016_ AuI._0017_ vssd1 vssd1 vccd1 vccd1 AuI._0018_ sky130_fd_sc_hd__and3_1
XANTENNA__10153__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07547__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._671_ AuI.pe._211_ AuI.pe._025_ AuI.pe._041_ AuI.pe._120_ AuI.pe._036_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._220_ sky130_fd_sc_hd__a221o_1
XANTENNA__07547__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A1 _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4742_ MuI._2852_ MuI._2884_ MuI._2880_ MuI.a_operand\[17\] vssd1 vssd1 vccd1
+ vccd1 MuI._0459_ sky130_fd_sc_hd__a22oi_1
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12540__B2 _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11169_ _06608_ _03051_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__nand2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1596_ AuI._0599_ vssd1 vssd1 vccd1 vccd1 AuI._0769_ sky130_fd_sc_hd__clkbuf_2
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08839__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4673_ MuI._0381_ MuI._0382_ vssd1 vssd1 vccd1 vccd1 MuI._0384_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5682__A2 MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6412_ MuI._2283_ MuI._2295_ vssd1 vssd1 vccd1 vccd1 MuI._2296_ sky130_fd_sc_hd__nor2_1
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3624_ MuI._1593_ MuI._1615_ vssd1 vssd1 vccd1 vccd1 MuI._2220_ sky130_fd_sc_hd__xor2_1
XANTENNA__07462__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6343_ MuI._2218_ MuI._2219_ vssd1 vssd1 vccd1 vccd1 MuI._2221_ sky130_fd_sc_hd__or2_1
XMuI._3555_ MuI.a_operand\[18\] vssd1 vssd1 vccd1 vccd1 MuI._1461_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5434__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__D _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ _06558_ _06571_ _06570_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__a21o_1
XMuI._6274_ MuI._2107_ MuI._2144_ vssd1 vssd1 vccd1 vccd1 MuI._2145_ sky130_fd_sc_hd__and2b_1
XMuI._3486_ MuI._0350_ MuI._0471_ MuI._0537_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._0702_
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13399__A3 _06306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08380_ _00993_ _00995_ _00994_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5225_ MuI._0947_ MuI._0950_ MuI._0989_ vssd1 vssd1 vccd1 vccd1 MuI._0991_ sky130_fd_sc_hd__and3_1
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07331_ _06630_ _06605_ _06591_ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a22oi_1
XFILLER_149_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5156_ MuI.a_operand\[14\] MuI.a_operand\[13\] MuI._0017_ MuI._0018_ vssd1 vssd1
+ vccd1 vccd1 MuI._0915_ sky130_fd_sc_hd__and4_1
XFILLER_137_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _06516_ _06562_ _06476_ _06520_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a22o_1
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4107_ MuI._2804_ MuI._2801_ vssd1 vssd1 vccd1 vccd1 MuI._3207_ sky130_fd_sc_hd__nor2_1
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _01616_ _01617_ _01611_ _01615_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a211o_1
XFILLER_118_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5087_ MuI._0836_ MuI._0832_ vssd1 vssd1 vccd1 vccd1 MuI._0839_ sky130_fd_sc_hd__xnor2_1
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07193_ net37 vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__buf_4
XFILLER_118_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4038_ MuI._3136_ MuI._3137_ vssd1 vssd1 vccd1 vccd1 MuI._3138_ sky130_fd_sc_hd__nor2_1
XFILLER_118_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06822__A _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12543__B _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3862__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _02556_ _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__nand2_1
XMuI._5989_ MuI._1795_ MuI._1814_ MuI._1808_ vssd1 vssd1 vccd1 vccd1 MuI._1831_ sky130_fd_sc_hd__a21o_1
XANTENNA__11159__B _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ _02404_ _02405_ _02487_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__or3_1
XANTENNA__12531__B2 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07653__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._515__A1 AuI.pe._070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09765_ _02411_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__xor2_1
X_06977_ _05176_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__buf_4
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08468__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11098__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _06500_ _04778_ _04832_ _06501_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__a22oi_2
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09696_ _02325_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__xnor2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09160__B1 _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _01166_ _01167_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__nor2_1
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13390__A _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ _01193_ _01187_ _01194_ _01195_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a211o_2
XFILLER_168_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _00144_ _00145_ _00069_ _00106_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__o211ai_2
XANTENNA__09299__B _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10073__A2 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _02431_ _02229_ _00163_ _03247_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__nand4_1
XANTENNA_MuI._3756__B MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _03170_ _03171_ _02989_ _02993_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__o211a_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12734__A _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _05043_ _05044_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ _02841_ _02910_ _02838_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a21o_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06732__A _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3772__A MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12141_ _04968_ _04969_ _04958_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3491__B MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12072_ _04736_ _02765_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__or2b_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11023_ _03764_ _03765_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__and3_1
XFILLER_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1450_ AuI._0422_ AuI._0424_ AuI._0428_ vssd1 vssd1 vccd1 vccd1 AuI._0636_ sky130_fd_sc_hd__and3_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._506__A1 AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1381_ AuI._0534_ AuI._0570_ AuI._0571_ AuI._0572_ vssd1 vssd1 vccd1 vccd1 AuI._0573_
+ sky130_fd_sc_hd__a211o_2
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10701__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12974_ _05797_ _05798_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__or2_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12286__B1 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6307__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__B1 _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _04722_ _04587_ _04738_ _04739_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__a211o_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4624__B1 MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _02905_ _02959_ _03449_ _05767_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__nand4_1
XFILLER_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06907__A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12628__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _03532_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__xnor2_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ _04570_ _04589_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__nand3_2
XANTENNA__09454__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5010_ MuI._0753_ vssd1 vssd1 vccd1 vccd1 MuI._0754_ sky130_fd_sc_hd__inv_2
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09454__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6377__B1 MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _03458_ _03459_ _03446_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a21o_1
XFILLER_159_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0856__A2 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13457_ _01322_ _01327_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2_1
XFILLER_174_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10669_ _03381_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__nand3_1
XANTENNA__08841__B _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0897__B AuI._0116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _05244_ _05245_ _05248_ _03315_ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__a221o_1
XANTENNA__11013__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11013__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13388_ _05883_ _06258_ _02817_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__a21bo_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12363__B _05047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5912_ MuI._1743_ MuI._1744_ MuI._1745_ vssd1 vssd1 vccd1 vccd1 MuI._1746_ sky130_fd_sc_hd__a21o_1
XFILLER_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12339_ _05061_ _05062_ _05064_ _05065_ _05056_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__a32o_1
XFILLER_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__A _02765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__B1 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5843_ MuI._1606_ MuI._1605_ vssd1 vssd1 vccd1 vccd1 MuI._1671_ sky130_fd_sc_hd__or2b_1
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13305__A3 _06209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._723_ AuI.pe._259_ AuI.pe._260_ AuI.pe._267_ AuI.pe._268_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._269_ sky130_fd_sc_hd__or4_1
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06900_ net34 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__buf_4
XMuI._5774_ MuI._1591_ MuI._1592_ MuI._1594_ vssd1 vssd1 vccd1 vccd1 MuI._1595_ sky130_fd_sc_hd__and3_1
XFILLER_141_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1648_ AuI.exp_a AuI.operand_a\[24\] AuI._0710_ AuI.operand_a\[25\] vssd1 vssd1
+ vccd1 vccd1 AuI._0004_ sky130_fd_sc_hd__a31o_1
X_07880_ _00495_ _00496_ _00350_ _00353_ vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__o211a_1
XFILLER_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._654_ AuI.pe._170_ AuI.pe._041_ AuI.pe._096_ AuI.pe._393_ AuI.pe._203_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._204_ sky130_fd_sc_hd__a221o_1
XFILLER_122_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4725_ MuI._0437_ MuI._0429_ MuI._0436_ vssd1 vssd1 vccd1 vccd1 MuI._0441_ sky130_fd_sc_hd__nand3_1
X_06831_ _03604_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11707__B _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1579_ AuI._0736_ AuI._0753_ AuI._0643_ vssd1 vssd1 vccd1 vccd1 AuI._0754_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._585_ AuI.pe._373_ AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 AuI.pe._140_ sky130_fd_sc_hd__or2_1
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4656_ MuI._0226_ MuI._0227_ MuI._0252_ vssd1 vssd1 vccd1 vccd1 MuI._0365_ sky130_fd_sc_hd__o21a_1
X_09550_ _02174_ _02176_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__and2_1
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06762_ _02862_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__and3_1
XMuI._3607_ MuI._0383_ MuI._0625_ MuI._1043_ MuI._1494_ vssd1 vssd1 vccd1 vccd1 MuI._2033_
+ sky130_fd_sc_hd__and4_1
XANTENNA__10330__C _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08501_ _01066_ _01067_ _01117_ _01118_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__nand4_1
XMuI._4587_ MuI._0286_ MuI._0287_ MuI._0288_ vssd1 vssd1 vccd1 vccd1 MuI._0289_ sky130_fd_sc_hd__o21ba_1
X_09481_ _01975_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or3_1
X_06693_ net2 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__clkinv_2
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12819__A _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6326_ MuI._2188_ MuI._2189_ vssd1 vssd1 vccd1 vccd1 MuI._2202_ sky130_fd_sc_hd__nor2_1
XFILLER_64_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3538_ MuI._1263_ vssd1 vssd1 vccd1 vccd1 MuI._1274_ sky130_fd_sc_hd__clkbuf_4
X_08432_ _01017_ _01018_ _01048_ _01049_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__and4bb_1
XFILLER_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06817__A _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6257_ MuI._2119_ MuI._2125_ vssd1 vssd1 vccd1 vccd1 MuI._2126_ sky130_fd_sc_hd__xnor2_1
XMuI._3469_ MuI._0504_ vssd1 vssd1 vccd1 vccd1 MuI._0515_ sky130_fd_sc_hd__clkbuf_4
X_08363_ _00979_ _00980_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__nor2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5208_ MuI._0969_ MuI._0970_ MuI._0971_ vssd1 vssd1 vccd1 vccd1 MuI._0972_ sky130_fd_sc_hd__nand3_1
XANTENNA__12257__C _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ _06609_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__nor2_1
XFILLER_177_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6188_ MuI._2046_ MuI._2049_ vssd1 vssd1 vccd1 vccd1 MuI._2050_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11252__B2 _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _03293_ _04046_ _04122_ _03239_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__a22o_1
XMuI._5139_ MuI._0866_ MuI._0870_ MuI._0868_ vssd1 vssd1 vccd1 vccd1 MuI._0896_ sky130_fd_sc_hd__o21ba_1
XFILLER_109_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07245_ _06489_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__buf_4
XFILLER_192_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07648__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__buf_4
XANTENNA__09566__C _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1415__C AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10763__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5894__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08479__A _00923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09817_ _02455_ _02456_ _02442_ _03884_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__o211a_1
XANTENNA__11617__B _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ _02347_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__or2_1
XFILLER_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07533__D net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _02320_ _02267_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__nor2_1
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09684__A1 _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__A _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11710_ _02723_ _05970_ _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__and3_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _05435_ _05491_ _05559_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__o211ai_2
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06727__A _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3767__A MuI._2866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11641_ _00445_ _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11243__A1 _03692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _04310_ _04324_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__nand2_1
XFILLER_168_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1309__D AuI._0506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _02830_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__or2_1
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 a_operand[22] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_6
X_10523_ _06593_ _05445_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__and2_1
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0950_ AuI._0110_ AuI._0157_ AuI._0159_ AuI._0161_ vssd1 vssd1 vccd1 vccd1 AuI._0162_
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _06150_ _06082_ _02837_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _03153_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__nor2_2
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0881_ net21 net113 vssd1 vssd1 vccd1 vccd1 AuI._0101_ sky130_fd_sc_hd__xor2_1
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11546__A2 _02931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12743__A1 _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _04211_ _04677_ _06079_ _06076_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__a211o_1
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10385_ net28 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__buf_2
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _04823_ _04824_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a21oi_2
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4748__D MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4763__A2_N MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1502_ AuI._0583_ AuI._0586_ vssd1 vssd1 vccd1 vccd1 AuI._0688_ sky130_fd_sc_hd__and2_1
XFILLER_105_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12055_ _04872_ _04878_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._3896__A1 MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3896__B2 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _03746_ _03747_ _03742_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__a21o_1
XAuI._1433_ AuI._0614_ AuI._0618_ vssd1 vssd1 vccd1 vccd1 AuI._0619_ sky130_fd_sc_hd__nand2_1
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10431__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4510_ MuI._0202_ MuI._0203_ vssd1 vssd1 vccd1 vccd1 MuI._0204_ sky130_fd_sc_hd__and2_1
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5490_ MuI._1272_ MuI._1280_ MuI._1227_ MuI._1281_ vssd1 vssd1 vccd1 vccd1 MuI._1282_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1364_ AuI._0438_ AuI._0333_ AuI._0498_ vssd1 vssd1 vccd1 vccd1 AuI._0557_ sky130_fd_sc_hd__or3_2
XANTENNA__07443__D _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4441_ MuI._0077_ MuI._0126_ MuI._0127_ vssd1 vssd1 vccd1 vccd1 MuI._0128_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _02809_ _05846_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__nand2_1
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1295_ AuI._0437_ AuI._0491_ AuI._0492_ AuI._0493_ vssd1 vssd1 vccd1 vccd1 AuI._0494_
+ sky130_fd_sc_hd__and4_1
XFuI._133__139 vssd1 vssd1 vccd1 vccd1 FuI._133__139/HI net139 sky130_fd_sc_hd__conb_1
XFILLER_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4372_ MuI._2440_ MuI._2975_ MuI._2976_ MuI._2671_ vssd1 vssd1 vccd1 vccd1 MuI._0053_
+ sky130_fd_sc_hd__a22oi_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _04719_ _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__xnor2_2
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6111_ MuI._0339_ MuI._2851_ MuI._2975_ MuI._0515_ vssd1 vssd1 vccd1 vccd1 MuI._1965_
+ sky130_fd_sc_hd__a22oi_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09383__A2_N _04111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12888_ _05772_ _02906_ _04635_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__mux2_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__A2 _03906_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5270__B1 MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _04736_ _02719_ _02722_ _02723_ _04645_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__a221o_1
XFILLER_187_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6042_ MuI._1887_ MuI._1888_ vssd1 vssd1 vccd1 vccd1 MuI._1889_ sky130_fd_sc_hd__xor2_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5022__B1 MuI._0725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__B1 _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ net25 vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07468__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12093__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI.pe._595__A AuI.pe._378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6875_ MuI._2501_ MuI._0174_ vssd1 vssd1 vccd1 vccd1 MuI._2775_ sky130_fd_sc_hd__and2b_1
XFILLER_142_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _02377_ _04714_ _01333_ _01334_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5826_ MuI._1164_ MuI._0421_ vssd1 vssd1 vccd1 vccd1 MuI._1652_ sky130_fd_sc_hd__nand2_1
XFILLER_142_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07932_ _04896_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__buf_4
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._706_ AuI.pe._072_ AuI.pe._164_ AuI.pe._225_ AuI.pe._013_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._253_ sky130_fd_sc_hd__a22o_1
XANTENNA__08166__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4955__B MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5757_ MuI._2836_ MuI._2838_ MuI._3349_ MuI._0085_ vssd1 vssd1 vccd1 vccd1 MuI._1576_
+ sky130_fd_sc_hd__nand4_1
XFILLER_69_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07863_ _00479_ _00478_ _00371_ _00212_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__o211ai_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6228__A MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._637_ AuI.pe._105_ AuI.pe._078_ AuI.pe._097_ AuI.pe._089_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._188_ sky130_fd_sc_hd__a22o_1
XFILLER_110_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07913__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4708_ MuI._0421_ MuI._0471_ MuI._0318_ MuI._0316_ MuI._0112_ vssd1 vssd1 vccd1
+ vccd1 MuI._0422_ sky130_fd_sc_hd__a32o_1
XFILLER_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5132__A MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ _02202_ _02193_ _02201_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nand3_1
XANTENNA__07913__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ net54 vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5688_ MuI._1482_ MuI._1498_ MuI._1499_ vssd1 vssd1 vccd1 vccd1 MuI._1500_ sky130_fd_sc_hd__nand3_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4836__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07794_ _05305_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__buf_4
XAuI.pe._568_ AuI.pe._046_ AuI.pe._086_ AuI.pe._123_ vssd1 vssd1 vccd1 vccd1 AuI.pe._124_
+ sky130_fd_sc_hd__a21o_1
XMuI._4639_ MuI._0343_ MuI._0345_ vssd1 vssd1 vccd1 vccd1 MuI._0346_ sky130_fd_sc_hd__nor2_1
X_09533_ _02090_ _02161_ _02163_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and3_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06745_ _02669_ _02615_ _02680_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__and3_1
XAuI.pe._499_ AuI.pe._059_ AuI.pe._049_ AuI.pe._060_ vssd1 vssd1 vccd1 vccd1 AuI.pe._061_
+ sky130_fd_sc_hd__o21a_1
X_09464_ _02074_ _02087_ _02069_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07650__B _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6309_ MuI._2178_ MuI._2182_ vssd1 vssd1 vccd1 vccd1 MuI._2183_ sky130_fd_sc_hd__xor2_2
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08415_ _01029_ _01032_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__xnor2_2
XFILLER_169_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11172__B _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09395_ _02009_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nand3_1
XFILLER_178_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ _00957_ _00962_ _00961_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a21o_1
XFILLER_132_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08277_ _00599_ _00598_ _00590_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__and2b_1
XFILLER_137_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07159_ net111 vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4211__A MuI._1021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09593__A _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _05058_ _03024_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__or2b_1
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout130 net24 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08157__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08157__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10889__D _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6138__A MuI._1993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07841__A _03324_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _01147_ _05948_ _05689_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__and3_1
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09657__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12459__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _00290_ _00289_ _03425_ _00163_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__nand4_1
XAuI._1080_ AuI._0180_ AuI._0187_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0291_ sky130_fd_sc_hd__mux2_1
XFILLER_188_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B1 _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08375__C net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _05540_ _05541_ _05451_ _05453_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o211ai_1
XANTENNA_MuI._5252__B1 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11624_ _04414_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__and2b_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09768__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12964__A1 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ _04339_ _04340_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o21a_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10707__A _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ _03209_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__or2b_1
XANTENNA__07288__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0933_ net21 AuI._0119_ AuI._0120_ vssd1 vssd1 vccd1 vccd1 AuI._0145_ sky130_fd_sc_hd__or3_1
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__xor2_4
XFILLER_183_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13225_ _06130_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__xnor2_1
XMuI._4990_ MuI._0730_ MuI._0731_ vssd1 vssd1 vccd1 vccd1 MuI._0732_ sky130_fd_sc_hd__or2_1
X_10437_ _02957_ _03003_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__o21ai_4
XAuI._0864_ AuI._0080_ net106 AuI._0082_ net36 vssd1 vssd1 vccd1 vccd1 AuI._0084_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10161__A_N _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3941_ MuI._0559_ MuI._0768_ MuI._2853_ MuI._2854_ vssd1 vssd1 vccd1 vccd1 MuI._3041_
+ sky130_fd_sc_hd__and4_1
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ _06058_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_2
X_10368_ _03044_ _03061_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__and3_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6747__S MuI._2487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06920__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6660_ MuI._0782_ MuI._2507_ vssd1 vssd1 vccd1 vccd1 MuI._2569_ sky130_fd_sc_hd__nor2_1
X_12107_ _04917_ _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__xor2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._1352__A AuI._0498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3872_ MuI._2969_ MuI._2970_ MuI._2971_ vssd1 vssd1 vccd1 vccd1 MuI._2972_ sky130_fd_sc_hd__a21bo_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _05938_ _05939_ _05985_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__a21oi_1
X_10299_ _02979_ _02986_ _02988_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__nand3_2
XMuI._5611_ MuI._3403_ MuI._0112_ MuI._1414_ vssd1 vssd1 vccd1 vccd1 MuI._1415_ sky130_fd_sc_hd__and3_1
XANTENNA__07139__A2_N _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6591_ MuI._0306_ MuI._2491_ MuI._2492_ vssd1 vssd1 vccd1 vccd1 MuI._2493_ sky130_fd_sc_hd__a21o_1
X_12038_ _04858_ _04859_ _04702_ _04749_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o211a_1
XFILLER_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10161__B _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5542_ MuI._1336_ MuI._1337_ MuI._1338_ vssd1 vssd1 vccd1 vccd1 MuI._1339_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4494__C MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1416_ AuI._0602_ vssd1 vssd1 vccd1 vccd1 AuI._0603_ sky130_fd_sc_hd__inv_2
XFILLER_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._422_ AuI.pe.significand\[13\] AuI.pe.significand\[14\] AuI.pe.significand\[15\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._389_ sky130_fd_sc_hd__nor3_1
XFILLER_207_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5473_ MuI._1207_ MuI._1262_ vssd1 vssd1 vccd1 vccd1 MuI._1264_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5887__A MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1347_ net13 net119 AuI._0126_ vssd1 vssd1 vccd1 vccd1 AuI._0542_ sky130_fd_sc_hd__mux2_2
XFILLER_207_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5102__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4424_ MuI.a_operand\[2\] vssd1 vssd1 vccd1 vccd1 MuI._0110_ sky130_fd_sc_hd__buf_2
XANTENNA__11273__A _02712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11704__C _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1278_ AuI._0476_ AuI._0477_ vssd1 vssd1 vccd1 vccd1 AuI._0478_ sky130_fd_sc_hd__xor2_4
XFILLER_209_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4355_ MuI._0027_ MuI._0033_ MuI._0034_ vssd1 vssd1 vccd1 vccd1 MuI._0035_ sky130_fd_sc_hd__a21oi_2
XFILLER_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3838__C MuI._2484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08200_ _00664_ _00663_ _06458_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a21o_1
XMuI._4286_ MuI._3383_ MuI._3385_ vssd1 vssd1 vccd1 vccd1 MuI._3386_ sky130_fd_sc_hd__or2b_1
X_09180_ _01784_ _01796_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__o21a_1
XFILLER_187_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6025_ MuI._3105_ MuI._1863_ MuI._1869_ vssd1 vssd1 vccd1 vccd1 MuI._1871_ sky130_fd_sc_hd__nor3_1
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12955__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _00713_ _00748_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__xor2_2
XFILLER_147_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07198__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08062_ _00677_ _00679_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__nor2_1
XANTENNA__10430__A2 _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07629__C _00246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6230__B MuI._0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10336__B _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07013_ _05563_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4669__C MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout106_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6858_ MuI._2735_ MuI._2760_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[23\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__11448__A _02593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08964_ _01580_ _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5809_ MuI._1573_ MuI._1631_ MuI._1632_ vssd1 vssd1 vccd1 vccd1 MuI._1633_ sky130_fd_sc_hd__and3_1
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6789_ MuI.Exception MuI._2710_ vssd1 vssd1 vccd1 vccd1 MuI._2711_ sky130_fd_sc_hd__and2b_1
XFILLER_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11167__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _00529_ _00531_ _00532_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__o21ba_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _01472_ _01479_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__nand2_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11694__A1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _00095_ _00096_ _04703_ _06611_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__and4_1
XANTENNA__08757__A _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07661__A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07777_ _00160_ _00165_ _00161_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__o21bai_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08476__B _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06728_ _02496_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__and3_1
X_09516_ _01981_ _01991_ _01990_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07380__B _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4037__A1 MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _06630_ net115 _03960_ _06631_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a22oi_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4037__B2 MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09588__A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _01981_ _01992_ _01993_ _01994_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a211o_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._102_ FuI._052_ FuI._060_ FuI.a_operand\[10\] vssd1 vssd1 vccd1 vccd1 FuI._000_
+ sky130_fd_sc_hd__o21a_1
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3467__D MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ _00908_ _00944_ _00945_ _00946_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__a211oi_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09811__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11340_ _03871_ _03872_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10421__A2 _00812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _02658_ _00783_ _05884_ _02593_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a22oi_2
XFILLER_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12742__A _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ _05782_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__nand2_1
XFILLER_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10222_ _02904_ _02804_ _02803_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a21o_1
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12461__B _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _03507_ _05671_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and2_1
XFILLER_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _01988_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__nand2_2
XANTENNA_input36_A a_operand[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12888__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09770__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07889__B1 _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12882__B1 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07571__A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1201_ AuI._0330_ AuI._0336_ AuI._0337_ AuI._0153_ vssd1 vssd1 vccd1 vccd1 AuI._0406_
+ sky130_fd_sc_hd__o31a_1
XFILLER_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11093__A _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11437__A1 _04076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1132_ AuI._0263_ AuI._0335_ AuI._0340_ AuI._0246_ vssd1 vssd1 vccd1 vccd1 AuI._0341_
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10986_ _03715_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4761__D MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _05522_ _05524_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__or2_1
XAuI._1063_ AuI._0206_ vssd1 vssd1 vccd1 vccd1 AuI._0274_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._4116__A MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12917__A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4140_ MuI._3237_ MuI._3239_ vssd1 vssd1 vccd1 vccd1 MuI._3240_ sky130_fd_sc_hd__nor2_1
XFILLER_204_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12656_ _05522_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06915__A _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__B _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4071_ MuI._3168_ MuI._3169_ MuI._3170_ vssd1 vssd1 vccd1 vccd1 MuI._3171_ sky130_fd_sc_hd__a21oi_2
XANTENNA_MuI._3955__A MuI._0581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08833__C _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ _04195_ _04194_ _04193_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__a21bo_1
X_12587_ _05446_ _05449_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__nand3_2
XANTENNA__09802__A1 _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09802__B2 _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _04312_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or2b_1
XFILLER_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0916_ AuI._0133_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[25\] sky130_fd_sc_hd__buf_2
X_11469_ _04222_ _04223_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__a21oi_2
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4973_ MuI._0710_ MuI._0712_ vssd1 vssd1 vccd1 vccd1 MuI._0714_ sky130_fd_sc_hd__nor2_1
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _06112_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__xor2_1
XAuI._0847_ net120 vssd1 vssd1 vccd1 vccd1 AuI._0067_ sky130_fd_sc_hd__inv_2
XFILLER_152_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6712_ MuI._2622_ MuI._2625_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2626_ sky130_fd_sc_hd__mux2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3924_ MuI._3022_ MuI._3023_ vssd1 vssd1 vccd1 vccd1 MuI._3024_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11912__A2 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _05947_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__inv_2
XFILLER_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6643_ MuI._1443_ MuI._2545_ MuI._2546_ MuI._2549_ vssd1 vssd1 vccd1 vccd1 MuI._2551_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_140_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3855_ MuI._2835_ MuI._2953_ MuI._2954_ vssd1 vssd1 vccd1 vccd1 MuI._2955_ sky130_fd_sc_hd__a21o_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._139__145 vssd1 vssd1 vccd1 vccd1 FuI._139__145/HI net145 sky130_fd_sc_hd__conb_1
X_07700_ _00092_ _00101_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__and2b_1
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6574_ MuI._2467_ MuI._2471_ MuI._2474_ vssd1 vssd1 vccd1 vccd1 MuI._2475_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13483__A _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3786_ MuI._2885_ vssd1 vssd1 vccd1 vccd1 MuI._2886_ sky130_fd_sc_hd__buf_2
XFILLER_94_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10479__A2 _03046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ _01291_ _01295_ _01296_ _01297_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__a211oi_4
XANTENNA_MuI._5113__C MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__B1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5525_ MuI._1260_ MuI._1267_ MuI._1268_ vssd1 vssd1 vccd1 vccd1 MuI._1321_ sky130_fd_sc_hd__and3_1
XANTENNA__07344__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07631_ _00020_ _00021_ _00247_ _00248_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__a211o_1
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08541__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._405_ AuI.pe._371_ vssd1 vssd1 vccd1 vccd1 AuI.pe._372_ sky130_fd_sc_hd__buf_2
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5464__B1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5456_ MuI._2881_ MuI._3245_ MuI._0304_ MuI._2892_ vssd1 vssd1 vccd1 vccd1 MuI._1245_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07562_ _00174_ _00178_ _00179_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__and3_1
XFILLER_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4407_ MuI._0081_ MuI._0083_ vssd1 vssd1 vccd1 vccd1 MuI._0091_ sky130_fd_sc_hd__xnor2_1
X_09301_ _02916_ _03917_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__and3_1
XMuI._5387_ MuI._1158_ MuI._1159_ vssd1 vssd1 vccd1 vccd1 MuI._1169_ sky130_fd_sc_hd__nand2_1
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07493_ _02948_ _04778_ _06603_ _02894_ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4026__A MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3568__C MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4338_ MuI._3388_ MuI._0004_ vssd1 vssd1 vccd1 vccd1 MuI._0016_ sky130_fd_sc_hd__xnor2_1
X_09232_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__or2_1
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12546__B _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__C _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4269_ MuI._0361_ MuI._0614_ MuI._2830_ MuI._3247_ vssd1 vssd1 vccd1 vccd1 MuI._3369_
+ sky130_fd_sc_hd__and4_1
X_09163_ _01772_ _01774_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6241__A MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6008_ MuI._3135_ MuI._3137_ MuI._3136_ vssd1 vssd1 vccd1 vccd1 MuI._1852_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10939__B1 _02707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5519__A1 MuI._2967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08114_ _00077_ _04531_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__nand2_1
XFILLER_135_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11600__A1 _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09094_ _06680_ _04305_ _01366_ _01367_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ _00527_ _00528_ _00661_ _00662_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__a211o_2
XANTENNA__12562__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13353__B2 _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3950__B1 MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _01316_ _01315_ _01275_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13105__A1 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13105__B2 _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08780__A1 _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4846__D MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08780__B2 _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _01547_ _01548_ _01562_ _01563_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__or4bb_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13393__A _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _01492_ _01494_ _01493_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a21o_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07391__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07829_ _00063_ _00216_ _06605_ _06591_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__nand4_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _03388_ _03387_ _03386_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a21bo_1
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08637__D _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10890__A2 _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _04197_ _02717_ _02730_ AuI.result\[3\] _03495_ vssd1 vssd1 vccd1 vccd1 _03496_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12092__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12092__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5758__A1 MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _02400_ _02584_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._5758__B2 MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ _06404_ _06358_ _06361_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nand3_1
XANTENNA__06735__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3775__A MuI._2868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ _05292_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__nor2_1
XFILLER_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09468__D net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ _05201_ _05202_ _05218_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o21ba_1
XFILLER_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ _04088_ _04089_ _03959_ _04054_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o211a_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ _02757_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__xor2_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10205_ _02442_ _04327_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__and2b_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ _03919_ _03941_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__and3_1
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3941__C MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__A1 _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _03842_ _05992_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__or2_1
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08771__B2 _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3640_ MuI.b_operand\[21\] MuI._2363_ MuI._2385_ MuI.b_operand\[22\] vssd1 vssd1
+ vccd1 vccd1 MuI._2396_ sky130_fd_sc_hd__a22o_1
XFILLER_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10067_ _02064_ _02020_ _06023_ _02705_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__and4b_1
XANTENNA__11658__A1 _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6238__A2 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3571_ MuI._1626_ MuI._0955_ vssd1 vssd1 vccd1 vccd1 MuI._1637_ sky130_fd_sc_hd__xnor2_1
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5310_ MuI._1067_ MuI._1083_ MuI._1081_ vssd1 vssd1 vccd1 vccd1 MuI._1084_ sky130_fd_sc_hd__a21o_1
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5230__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6290_ MuI._2126_ MuI._2139_ vssd1 vssd1 vccd1 vccd1 MuI._2162_ sky130_fd_sc_hd__nor2_1
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09079__A2 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5241_ MuI._1002_ MuI._1007_ vssd1 vssd1 vccd1 vccd1 MuI._1008_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1115_ AuI._0254_ AuI._0301_ AuI._0300_ vssd1 vssd1 vccd1 vccd1 AuI._0325_ sky130_fd_sc_hd__a21bo_1
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12720__A_N _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _03524_ _03526_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__and2_1
XFILLER_204_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08844__B _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5172_ MuI._2841_ MuI._0305_ vssd1 vssd1 vccd1 vccd1 MuI._0932_ sky130_fd_sc_hd__nand2_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1046_ AuI._0257_ vssd1 vssd1 vccd1 vccd1 AuI._0258_ sky130_fd_sc_hd__buf_2
X_12708_ _05363_ _02853_ _05373_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a31o_1
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4123_ MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 MuI._3223_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._3685__A MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4421__B2 MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4054_ MuI._3081_ MuI._3084_ MuI._3153_ vssd1 vssd1 vccd1 vccd1 MuI._3154_ sky130_fd_sc_hd__a21oi_2
XANTENNA__12085__C _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11697__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07262__A1 _06516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07262__B2 _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4956_ MuI._2837_ MuI.a_operand\[9\] MuI._2341_ MuI._2853_ vssd1 vssd1 vccd1
+ vccd1 MuI._0695_ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._4947__C MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _02502_ _02504_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__nand2_1
XFILLER_98_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07195__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11897__A1 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3907_ MuI._3004_ MuI._3005_ MuI._2996_ vssd1 vssd1 vccd1 vccd1 MuI._3007_ sky130_fd_sc_hd__a21oi_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08801_ _01416_ _01418_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nor2_2
XMuI._4887_ MuI._0616_ MuI._0618_ vssd1 vssd1 vccd1 vccd1 MuI._0619_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._4666__D MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _05349_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[21\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__13099__B1 _05998_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ _02428_ _02426_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__and2b_1
XFILLER_100_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10098__B_N _02496_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6626_ MuI._3397_ MuI._0421_ MuI._1436_ MuI._2531_ vssd1 vssd1 vccd1 vccd1 MuI._2532_
+ sky130_fd_sc_hd__a211o_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3838_ MuI.b_operand\[19\] MuI._2811_ MuI._2484_ MuI._2773_ vssd1 vssd1 vccd1
+ vccd1 MuI._2938_ sky130_fd_sc_hd__and4_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _00414_ _04509_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__nand2_2
XANTENNA_AuI.pe._542__A2 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09841__D _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6557_ MuI._2442_ MuI._2446_ MuI._2449_ MuI._2455_ vssd1 vssd1 vccd1 vccd1 MuI._2456_
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3769_ MuI._2868_ vssd1 vssd1 vccd1 vccd1 MuI._2869_ sky130_fd_sc_hd__clkbuf_4
XFILLER_94_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08738__C _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08663_ _06460_ _05101_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__nand2_1
XANTENNA__07642__C _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5508_ MuI._1300_ MuI._1301_ vssd1 vssd1 vccd1 vccd1 MuI._1302_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5140__A MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6488_ MuI._2378_ MuI._2379_ vssd1 vssd1 vccd1 vccd1 MuI._2380_ sky130_fd_sc_hd__nor2_1
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07614_ _00231_ _00083_ _00098_ _03217_ vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__a22o_1
XFILLER_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _01164_ _01168_ _01170_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__or3b_1
XFILLER_81_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5439_ MuI._1215_ MuI._1216_ MuI._1202_ MuI._1214_ vssd1 vssd1 vccd1 vccd1 MuI._1226_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ net130 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_MuI._6670__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11821__A1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _03163_ _00093_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__nand2_1
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11821__B2 _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09215_ _01784_ _01795_ _01789_ _01794_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__o211a_1
XFILLER_194_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1418__C AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__D _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09146_ _01761_ _01760_ _01758_ _01735_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__o211a_1
XFILLER_148_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08770__A _01382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ _01601_ _01598_ _01600_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__a21o_1
XFILLER_107_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ _00641_ _00644_ _00645_ _06641_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__o211ai_4
XFILLER_190_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12404__B1_N _06629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__B1 _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._781__A2 AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4479__A1 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4479__B2 MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _02633_ _02638_ _02642_ _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a211o_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10540__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._533__A2 AuI.pe._042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ _05809_ _05808_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or2b_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11941_ _04652_ _04653_ _04755_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a211oi_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4592__C MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12065__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _03548_ _03549_ _03363_ _03367_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__o211ai_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _03475_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__xnor2_2
XFILLER_201_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13473_ _02921_ _06338_ _02824_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__a21o_1
X_10685_ _03401_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21o_1
XFILLER_201_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09769__B1 _00266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _03099_ _00785_ _05884_ _03056_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a22oi_2
XFILLER_154_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6156__A1 MuI._0779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6156__B2 MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _05199_ _05200_ _05183_ _05107_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__o211a_1
XANTENNA__11040__A2 _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07795__A2 _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _00077_ _00197_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nand2_1
XFILLER_154_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12286_ _05033_ _05034_ _05126_ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__o211ai_2
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4810_ MuI._0456_ MuI._0533_ vssd1 vssd1 vccd1 vccd1 MuI._0534_ sky130_fd_sc_hd__xor2_2
XFILLER_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3914__B1 MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5790_ MuI._1609_ MuI._1610_ MuI._1611_ vssd1 vssd1 vccd1 vccd1 MuI._1612_ sky130_fd_sc_hd__nand3_1
XFILLER_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11237_ _03696_ _03823_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a21oi_4
XFILLER_84_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1664_ AuI.operand_a\[28\] AuI._0604_ AuI._0710_ vssd1 vssd1 vccd1 vccd1 AuI._0017_
+ sky130_fd_sc_hd__nand3_1
XFILLER_122_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12930__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._670_ AuI.pe._084_ AuI.pe._119_ AuI.pe._218_ AuI.pe._201_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._219_ sky130_fd_sc_hd__a22o_1
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4741_ MuI._2616_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._0458_ sky130_fd_sc_hd__nand2_1
XANTENNA__07547__A2 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12540__A2 _05702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11168_ _03922_ _03923_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__nor2_1
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1595_ AuI._0693_ AuI._0763_ AuI._0767_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0768_
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10551__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08839__B _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4672_ MuI._0150_ MuI._0149_ vssd1 vssd1 vccd1 vccd1 MuI._0382_ sky130_fd_sc_hd__and2b_1
X_10119_ _02792_ _02793_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__or2_1
X_11099_ _02545_ _02553_ _02565_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a21o_1
XFILLER_110_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10450__A _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6411_ MuI._2283_ MuI._2293_ MuI._2294_ vssd1 vssd1 vccd1 vccd1 MuI._2295_ sky130_fd_sc_hd__nor3_1
XFILLER_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3623_ MuI._2176_ MuI._2187_ MuI._2198_ vssd1 vssd1 vccd1 vccd1 MuI._2209_ sky130_fd_sc_hd__a21bo_1
XFILLER_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07462__C _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6342_ MuI._0372_ MuI._0625_ MuI._1494_ MuI._2077_ vssd1 vssd1 vccd1 vccd1 MuI._2219_
+ sky130_fd_sc_hd__and4_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3554_ MuI._1428_ MuI._1439_ vssd1 vssd1 vccd1 vccd1 MuI._1450_ sky130_fd_sc_hd__nor2_1
XFILLER_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6092__B1 MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6273_ MuI._2108_ MuI._2142_ vssd1 vssd1 vccd1 vccd1 MuI._2144_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3485_ MuI._0350_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._0691_ sky130_fd_sc_hd__nand2_1
XFILLER_91_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5224_ MuI._0947_ MuI._0950_ MuI._0989_ vssd1 vssd1 vccd1 vccd1 MuI._0990_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ _06598_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__buf_4
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11803__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5155_ MuI._0327_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0914_ sky130_fd_sc_hd__nand2_1
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07261_ net18 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__buf_4
XAuI._1029_ AuI._0239_ AuI._0240_ AuI._0223_ vssd1 vssd1 vccd1 vccd1 AuI._0241_ sky130_fd_sc_hd__mux2_1
XFILLER_176_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4106_ MuI._3204_ MuI._3201_ vssd1 vssd1 vccd1 vccd1 MuI._3206_ sky130_fd_sc_hd__xnor2_1
X_09000_ _01611_ _01615_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__o211ai_2
XFILLER_192_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6222__C MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5086_ MuI._2919_ MuI._0321_ vssd1 vssd1 vccd1 vccd1 MuI._0838_ sky130_fd_sc_hd__nand2_1
X_07192_ _06491_ _06466_ _06461_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__a22oi_2
XFILLER_157_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08590__A _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4037_ MuI._1494_ MuI._2800_ MuI._2919_ MuI._1032_ vssd1 vssd1 vccd1 vccd1 MuI._3137_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3862__B MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09902_ _02558_ _02560_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__and2_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5988_ MuI._1826_ MuI._1829_ vssd1 vssd1 vccd1 vccd1 MuI._1830_ sky130_fd_sc_hd__or2_1
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__C _03913_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4939_ MuI._2660_ MuI._2884_ MuI._3307_ MuI._2605_ vssd1 vssd1 vccd1 vccd1 MuI._0676_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_99_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09833_ _02449_ _02481_ _02441_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a21o_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._799_ AuI.operand_a\[25\] AuI.pe._331_ AuI.pe._333_ AuI.pe._338_ vssd1 vssd1
+ vccd1 vccd1 AuI.pe._339_ sky130_fd_sc_hd__and4_1
XFILLER_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09764_ _06475_ _03960_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__nand2_1
XANTENNA__10360__A _06593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06976_ net15 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__clkbuf_4
XMuI._6609_ MuI._1829_ MuI._2512_ vssd1 vssd1 vccd1 vccd1 MuI._2513_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08468__C _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08715_ _01332_ _02334_ _06611_ _06602_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__and4_1
XFILLER_55_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ _02336_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__or2_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09160__A1 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09160__B2 _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08646_ _01261_ _01252_ _01258_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__and3_1
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__A _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _00908_ _00941_ _00942_ _00943_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__and4_1
XFILLER_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07528_ _00069_ _00106_ _00144_ _00145_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__a211o_1
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09299__C _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07459_ net114 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._3756__C MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _02989_ _02993_ _03170_ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__a211oi_2
XFILLER_109_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12734__B _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09129_ _01737_ _01746_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__or2b_1
XFILLER_109_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1275__B1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._658__D AuI.pe._101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _04958_ _04968_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._3772__B MuI._2871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _03134_ _04879_ _04880_ _04891_ _04895_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a311o_4
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _03579_ _03581_ _03580_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__a21bo_1
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07844__A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4884__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._506__A2 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1380_ AuI._0555_ AuI._0561_ AuI._0562_ vssd1 vssd1 vccd1 vccd1 AuI._0572_ sky130_fd_sc_hd__a21boi_1
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10701__C _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12973_ _05784_ _05824_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and2_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09151__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09151__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _04735_ _04737_ _04579_ _04583_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__o211a_1
XANTENNA__10118__A_N _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _00216_ _05702_ _05767_ _00217_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._4624__B2 MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _03798_ _04262_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nand2_1
XFILLER_159_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11786_ _04587_ _04588_ _04460_ _04571_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a211o_1
XANTENNA__09454__A2 _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6377__A1 MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6377__B2 MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10737_ _03446_ _03458_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__nand3_2
XFILLER_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _02822_ _06369_ _02713_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06923__A _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10668_ _00221_ _05123_ _03382_ _03383_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nand4_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08841__C _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _05251_ _05254_ _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__or3_1
XANTENNA_AuI._1266__A0 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__A2 _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _03301_ _03305_ _03311_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__or3_1
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13387_ _06298_ _06300_ _06428_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__a21oi_1
XMuI._5911_ MuI._0701_ MuI._0704_ vssd1 vssd1 vccd1 vccd1 MuI._1745_ sky130_fd_sc_hd__xnor2_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07768__A2 _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ _05093_ _05103_ _05104_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nand3_1
XFILLER_181_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10164__B _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5842_ MuI._1598_ MuI._1603_ vssd1 vssd1 vccd1 vccd1 MuI._1669_ sky130_fd_sc_hd__or2b_1
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12269_ _04970_ _04973_ _05107_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o211ai_2
XFILLER_123_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._722_ AuI.pe._013_ AuI.pe._012_ AuI.pe._213_ AuI.pe._045_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._268_ sky130_fd_sc_hd__a22o_1
XFILLER_141_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5773_ MuI._1490_ MuI._1498_ vssd1 vssd1 vccd1 vccd1 MuI._1594_ sky130_fd_sc_hd__nand2_1
XAuI._1647_ AuI._0695_ AuI._0001_ AuI._0003_ vssd1 vssd1 vccd1 vccd1 AuI.result\[24\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._653_ AuI.pe.significand\[13\] AuI.pe._004_ AuI.pe._006_ AuI.pe._120_ AuI.pe._202_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._203_ sky130_fd_sc_hd__a221o_1
XFILLER_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4724_ MuI._0439_ vssd1 vssd1 vccd1 vccd1 MuI._0440_ sky130_fd_sc_hd__inv_2
XFILLER_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06830_ _03593_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__buf_2
XAuI._1578_ AuI._0638_ AuI._0639_ AuI._0667_ vssd1 vssd1 vccd1 vccd1 AuI._0753_ sky130_fd_sc_hd__and3_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._584_ AuI.pe._020_ AuI.pe._133_ AuI.pe._136_ AuI.pe._138_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._139_ sky130_fd_sc_hd__a211o_1
XMuI._4655_ MuI._0341_ MuI._0363_ MuI._0360_ vssd1 vssd1 vccd1 vccd1 MuI._0364_ sky130_fd_sc_hd__a21o_1
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06761_ _02851_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__buf_6
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4863__A1 MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4863__B2 MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3606_ MuI._0636_ MuI._1043_ MuI._1494_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._2022_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10330__D _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _01114_ _01115_ _01092_ _01105_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__o211ai_2
XMuI._4586_ MuI._2799_ MuI._2918_ MuI._3223_ MuI._3349_ vssd1 vssd1 vccd1 vccd1 MuI._0288_
+ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._5862__A1_N MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ _02101_ _02103_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a21bo_1
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06692_ _02107_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__buf_6
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08585__A _03239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6325_ MuI._2158_ MuI._2159_ vssd1 vssd1 vccd1 vccd1 MuI._2201_ sky130_fd_sc_hd__nand2_1
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3537_ MuI.b_operand\[17\] vssd1 vssd1 vccd1 vccd1 MuI._1263_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12819__B _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _01046_ _01047_ _01035_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a21o_1
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6256_ MuI._2123_ MuI._2124_ vssd1 vssd1 vccd1 vccd1 MuI._2125_ sky130_fd_sc_hd__xor2_1
XMuI._3468_ MuI._0482_ MuI._0493_ vssd1 vssd1 vccd1 vccd1 MuI._0504_ sky130_fd_sc_hd__nand2_1
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08362_ net110 net109 net14 _05176_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__and4_1
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5207_ MuI._0811_ MuI._0813_ vssd1 vssd1 vccd1 vccd1 MuI._0971_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11788__B1 _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07313_ _06610_ _06613_ _06600_ _06607_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_177_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6187_ MuI._2047_ MuI._2048_ vssd1 vssd1 vccd1 vccd1 MuI._2049_ sky130_fd_sc_hd__and2b_1
XANTENNA_AuI.pe._681__B2 AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__D _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _00608_ _00910_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__or2_1
XFILLER_177_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12835__A _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5138_ MuI._0883_ MuI._0884_ MuI._0894_ vssd1 vssd1 vccd1 vccd1 MuI._0895_ sky130_fd_sc_hd__nand3_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07244_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__buf_4
XFILLER_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06833__A _03626_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5069_ MuI._0815_ MuI._0818_ vssd1 vssd1 vccd1 vccd1 MuI._0819_ sky130_fd_sc_hd__xnor2_1
X_07175_ net19 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10355__A _03046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__D _00084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12570__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08479__B _00922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__inv_2
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09747_ _02393_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__inv_2
X_06959_ _04983_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__clkbuf_4
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ _02265_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__inv_2
XANTENNA__07144__B1 _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09684__A2 _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12729__B _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _06601_ _04445_ _00085_ _06606_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__a22oi_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _03604_ _06612_ _06603_ _06434_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a22o_1
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11571_ _04161_ _04350_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _06218_ _06219_ _02926_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__mux2_1
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _00000_ _02669_ _03051_ _03071_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__nand4_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06743__A _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3783__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13241_ _03400_ _05531_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__nand2_1
X_10453_ _03141_ _03142_ _03151_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__and3_1
XFILLER_109_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0880_ AuI._0098_ AuI._0099_ vssd1 vssd1 vccd1 vccd1 AuI._0100_ sky130_fd_sc_hd__nand2_2
XFILLER_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12743__A2 _03071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13172_ _03239_ _05338_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__nor2_1
XANTENNA_input66_A b_operand[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _06500_ _00785_ _00153_ _06501_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a22o_1
XFILLER_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12123_ _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__and2_1
XFILLER_151_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4542__B1 MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1501_ AuI._0596_ AuI._0598_ vssd1 vssd1 vccd1 vccd1 AuI._0687_ sky130_fd_sc_hd__and2_1
XFILLER_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12054_ _04872_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3896__A2 MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _03742_ _03746_ _03747_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nand3_1
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1432_ AuI._0389_ AuI._0449_ AuI._0422_ AuI._0550_ vssd1 vssd1 vccd1 vccd1 AuI._0618_
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07383__B1 _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1363_ AuI._0551_ AuI._0554_ AuI._0555_ vssd1 vssd1 vccd1 vccd1 AuI._0556_ sky130_fd_sc_hd__a21bo_1
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13456__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4440_ MuI._0075_ MuI._0076_ vssd1 vssd1 vccd1 vccd1 MuI._0127_ sky130_fd_sc_hd__nor2_1
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12956_ _02809_ _05846_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__or2_1
XFILLER_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1294_ net9 net41 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0493_ sky130_fd_sc_hd__mux2_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06918__A _04542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4371_ MuI._2850_ MuI._2539_ vssd1 vssd1 vccd1 vccd1 MuI._0052_ sky130_fd_sc_hd__nand2_1
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11907_ _03798_ _04736_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__nand2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6110_ MuI._1893_ MuI._1898_ vssd1 vssd1 vccd1 vccd1 MuI._1964_ sky130_fd_sc_hd__nand2_1
X_12887_ _02805_ _05685_ _02802_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__a21o_1
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _02723_ _04671_ _02744_ _04627_ FuI.Integer\[11\] vssd1 vssd1 vccd1 vccd1
+ _04645_ sky130_fd_sc_hd__a32o_1
XFILLER_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6041_ MuI.a_operand\[25\] MuI._2889_ MuI._2890_ MuI._2976_ vssd1 vssd1 vccd1
+ vccd1 MuI._1888_ sky130_fd_sc_hd__o31a_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ _04278_ _04282_ _04460_ _04461_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a211oi_2
XFILLER_159_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ _06332_ _06333_ _06341_ _02751_ _06353_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__a221o_4
XFILLER_174_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10175__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12093__C _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6874_ MuI._2735_ MuI._2774_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[28\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_103_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4870__A2_N MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08980_ _01592_ _01593_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a21o_1
XFILLER_170_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5825_ MuI._1574_ MuI._1589_ MuI._1590_ MuI._1595_ vssd1 vssd1 vccd1 vccd1 MuI._1651_
+ sky130_fd_sc_hd__a31o_1
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _00546_ _00548_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__nor2_1
XAuI.pe._705_ AuI.pe._142_ AuI.pe._097_ AuI.pe._246_ AuI.pe._251_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._252_ sky130_fd_sc_hd__a211o_1
XMuI._5756_ MuI.b_operand\[11\] MuI._3362_ vssd1 vssd1 vccd1 vccd1 MuI._1575_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._4955__C MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__A2 _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1411__B1 AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _00212_ _00371_ _00478_ _00479_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__a211o_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._636_ AuI.pe._059_ AuI.pe._133_ AuI.pe._173_ AuI.pe._029_ AuI.pe._186_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._187_ sky130_fd_sc_hd__a221o_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4707_ MuI._0420_ vssd1 vssd1 vccd1 vccd1 MuI._0421_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._6228__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _02226_ _02234_ _02236_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07913__A2 _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5132__B MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5687_ MuI._1490_ MuI._1491_ MuI._1497_ vssd1 vssd1 vccd1 vccd1 MuI._1499_ sky130_fd_sc_hd__a21o_1
X_06813_ _03411_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[24\] sky130_fd_sc_hd__clkbuf_1
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4029__A MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4836__A1 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07793_ _02712_ _06568_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__nand2_1
XFILLER_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4836__B2 MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4638_ MuI._0344_ MuI._0342_ vssd1 vssd1 vccd1 vccd1 MuI._0345_ sky130_fd_sc_hd__or2_1
XAuI.pe._567_ AuI.pe._063_ AuI.pe._066_ AuI.pe._054_ AuI.pe._072_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._123_ sky130_fd_sc_hd__a22o_1
XANTENNA__13425__S _04635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09532_ _02159_ _02160_ _02138_ _02143_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__o211ai_1
X_06744_ _02151_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__clkbuf_2
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._498_ AuI.pe._056_ AuI.pe._049_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._060_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_92_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4569_ MuI._0268_ MuI._0115_ vssd1 vssd1 vccd1 vccd1 MuI._0269_ sky130_fd_sc_hd__nor2_1
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _02081_ _02085_ _02074_ _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07650__C _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6308_ MuI._2180_ MuI._2181_ vssd1 vssd1 vccd1 vccd1 MuI._2182_ sky130_fd_sc_hd__xnor2_1
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _01030_ _01031_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and2b_1
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11172__C _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ _02009_ _02010_ _02011_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a21o_1
XANTENNA__10069__B _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6239_ MuI._2104_ MuI._2105_ vssd1 vssd1 vccd1 vccd1 MuI._2106_ sky130_fd_sc_hd__nor2_1
XFILLER_178_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._654__B2 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ _00957_ _00961_ _00962_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__nand3_1
XFILLER_177_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ _00599_ _00590_ _00598_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__and3_1
XFILLER_193_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__C _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07378__B _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ _06515_ net17 _05305_ _06519_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__a22o_1
XFILLER_165_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09874__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _02096_ _02194_ net23 net130 vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__and4_1
XANTENNA__09051__B1 _01668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4211__B MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07089_ _04865_ _06284_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__and2_1
XFILLER_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07394__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12489__A1 _05266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout120 net43 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
Xfanout131 net24 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08157__A2 _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _03239_ _05959_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07841__B _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09657__A2 _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12459__B _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _00279_ _00382_ _00163_ _03378_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a22o_1
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6154__A MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B2 _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08375__D net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5252__A1 MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12672_ _05451_ _05453_ _05540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a211o_1
XFILLER_169_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5252__B2 MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _04409_ _04410_ _04412_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__a21o_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09768__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11554_ _04339_ _04340_ _02713_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__a21oi_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10707__B _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ _03206_ _03207_ _03208_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a21o_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07288__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07840__A1 _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0932_ AuI._0128_ AuI._0129_ net53 vssd1 vssd1 vccd1 vccd1 AuI._0144_ sky130_fd_sc_hd__a21o_1
XFILLER_156_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _04105_ _04106_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a21oi_2
XANTENNA_MuI._4963__A1_N MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12177__B1 _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12716__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ _06047_ _06049_ _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a21o_1
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10436_ _03001_ _02958_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__or2b_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0863_ AuI._0078_ net6 AuI._0082_ net36 vssd1 vssd1 vccd1 vccd1 AuI._0083_ sky130_fd_sc_hd__o22ai_1
XMuI._3940_ MuI._1010_ MuI.b_operand\[11\] vssd1 vssd1 vccd1 vccd1 MuI._3040_ sky130_fd_sc_hd__nand2_1
XFILLER_98_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _05983_ _05984_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ _03059_ _03060_ _03050_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__a21o_1
XANTENNA__10723__A _02345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3871_ MuI._2968_ MuI._2964_ MuI._2965_ vssd1 vssd1 vccd1 vccd1 MuI._2971_ sky130_fd_sc_hd__nand3_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04923_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10298_ _02987_ _04380_ _02982_ _02985_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__nand4_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _05938_ _05939_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and3_1
XMuI._5610_ MuI._3397_ MuI._0245_ vssd1 vssd1 vccd1 vccd1 MuI._1414_ sky130_fd_sc_hd__and2_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10442__B _04133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6590_ MuI._0295_ MuI._0284_ MuI._0262_ vssd1 vssd1 vccd1 vccd1 MuI._2492_ sky130_fd_sc_hd__and3b_1
XFILLER_26_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12037_ _04702_ _04749_ _04858_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a211oi_1
XFILLER_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI.pe._581__B1 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5541_ MuI._2966_ MuI.a_operand\[0\] vssd1 vssd1 vccd1 vccd1 MuI._1338_ sky130_fd_sc_hd__and2_1
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1415_ AuI.exp_a AuI.operand_a\[24\] AuI.operand_a\[25\] vssd1 vssd1 vccd1 vccd1
+ AuI._0602_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._4494__D MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._421_ AuI.pe._382_ AuI.pe._384_ AuI.pe._387_ vssd1 vssd1 vccd1 vccd1 AuI.pe._388_
+ sky130_fd_sc_hd__and3_2
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5472_ MuI._1210_ MuI._1209_ vssd1 vssd1 vccd1 vccd1 MuI._1262_ sky130_fd_sc_hd__nor2_1
XAuI._1346_ AuI._0539_ AuI._0540_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0541_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._5887__B MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07293__A2_N _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4423_ MuI._0106_ MuI._0107_ vssd1 vssd1 vccd1 vccd1 MuI._0109_ sky130_fd_sc_hd__nor2_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12369__B _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3688__A MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11273__B _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _05826_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__and2_1
XAuI._1277_ net8 net40 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0477_ sky130_fd_sc_hd__mux2_4
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4354_ MuI._0024_ MuI._0026_ vssd1 vssd1 vccd1 vccd1 MuI._0034_ sky130_fd_sc_hd__and2_1
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._3838__D MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4285_ MuI._3382_ MuI._3384_ vssd1 vssd1 vccd1 vccd1 MuI._3385_ sky130_fd_sc_hd__and2_1
XFILLER_159_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6024_ MuI._3105_ MuI._1863_ MuI._1869_ vssd1 vssd1 vccd1 vccd1 MuI._1870_ sky130_fd_sc_hd__o21a_1
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _00746_ _00747_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__nand2_1
XFILLER_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07479__A _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _03539_ _00678_ _00287_ _00267_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__and4_1
XFILLER_174_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07198__B _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07012_ net22 vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12168__B1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12707__A2 _03186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4669__D MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09536__A1_N _06620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__A _00124_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6857_ MuI._2503_ MuI._2733_ MuI._2731_ MuI.Exception vssd1 vssd1 vccd1 vccd1
+ MuI._2761_ sky130_fd_sc_hd__a211o_2
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _01405_ _01407_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nor2_1
XANTENNA__11448__B _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5808_ MuI._1629_ MuI._1630_ MuI._1541_ MuI._1543_ vssd1 vssd1 vccd1 vccd1 MuI._1632_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ _06501_ _06500_ _06562_ _05370_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__and4_1
XMuI._6788_ MuI._2708_ MuI._2709_ vssd1 vssd1 vccd1 vccd1 MuI._2710_ sky130_fd_sc_hd__xnor2_1
XANTENNA_AuI.pe._572__B1 AuI.pe._079_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__C _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ _01473_ _01478_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__or2b_1
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5739_ MuI._1464_ MuI._1552_ MuI._1553_ vssd1 vssd1 vccd1 vccd1 MuI._1556_ sky130_fd_sc_hd__or3_1
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _00462_ _04703_ _04778_ _00237_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__a22oi_2
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._619_ AuI.pe._170_ AuI.pe._167_ vssd1 vssd1 vccd1 vccd1 AuI.pe._171_ sky130_fd_sc_hd__xor2_1
XANTENNA__08757__B _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _00177_ _00178_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__nand2_1
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _02127_ _02128_ _02135_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__nand3_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06727_ _02485_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__clkbuf_8
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ _02754_ _02797_ net115 net132 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__and4_2
XANTENNA_MuI._4037__A2 MuI._2800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._101_ FuI._037_ FuI._055_ vssd1 vssd1 vccd1 vccd1 FuI._060_ sky130_fd_sc_hd__and2_1
X_09377_ _01981_ _01992_ _01993_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09588__B _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11403__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08328_ _00653_ _00654_ _00620_ _00655_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__and4_1
XANTENNA__08075__A1 _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1437__B AuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__B2 _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09811__A2 _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._5318__A MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08259_ _06598_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__buf_4
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _04031_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12742__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _02867_ _02903_ _02866_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__o21ba_1
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _02828_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or2_2
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5053__A MuI._3189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10083_ _02442_ _04327_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__or2_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09770__C net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A a_operand[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1200_ AuI._0268_ AuI._0271_ AuI._0274_ vssd1 vssd1 vccd1 vccd1 AuI._0405_ sky130_fd_sc_hd__mux2_1
XANTENNA__07571__B _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1131_ AuI._0233_ AuI._0336_ AuI._0337_ AuI._0339_ AuI._0153_ vssd1 vssd1 vccd1
+ vccd1 AuI._0340_ sky130_fd_sc_hd__o311a_1
XANTENNA__11093__B _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _03724_ _03721_ _03723_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nand3_2
XFILLER_43_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12724_ _02868_ _05596_ _05597_ _02750_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__o211a_1
XAuI._1062_ AuI._0173_ AuI._0272_ AuI._0176_ vssd1 vssd1 vccd1 vccd1 AuI._0273_ sky130_fd_sc_hd__mux2_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4116__B MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12917__B _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12655_ _05431_ _05432_ _05523_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4070_ MuI._3165_ MuI._3167_ vssd1 vssd1 vccd1 vccd1 MuI._3170_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._3787__A1 MuI._0482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ _04394_ _04392_ _04393_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__nand3_1
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07299__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__C _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3955__B MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__D _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _03486_ _05456_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__nand4_2
XANTENNA__09802__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ _02703_ _04315_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__a21oi_2
XFILLER_156_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output97_A net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0915_ net22 net54 AuI._0121_ vssd1 vssd1 vccd1 vccd1 AuI._0133_ sky130_fd_sc_hd__mux2_1
XFILLER_144_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11468_ _04050_ _04246_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__xor2_1
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12652__B _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08591__A2_N _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4972_ MuI._0710_ MuI._0711_ MuI.b_operand\[14\] MuI._3246_ vssd1 vssd1 vccd1
+ vccd1 MuI._0712_ sky130_fd_sc_hd__and4bb_1
X_13207_ _03680_ _05713_ _06018_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a31o_1
X_10419_ _02952_ _03117_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__xnor2_1
XAuI._0846_ AuI._0061_ AuI._0063_ AuI._0065_ AuI._0052_ AuI._0055_ vssd1 vssd1 vccd1
+ vccd1 AuI._0066_ sky130_fd_sc_hd__a2111o_1
X_11399_ _04157_ _04160_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__a21oi_2
XMuI._6711_ MuI._2339_ MuI._2624_ vssd1 vssd1 vccd1 vccd1 MuI._2625_ sky130_fd_sc_hd__xnor2_1
XMuI._3923_ MuI._2385_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._3023_ sky130_fd_sc_hd__nand2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _06039_ _06040_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2_1
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1090__A1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6642_ MuI._1181_ MuI._2548_ vssd1 vssd1 vccd1 vccd1 MuI._2549_ sky130_fd_sc_hd__xnor2_1
XMuI._3854_ MuI._2926_ MuI._2952_ vssd1 vssd1 vccd1 vccd1 MuI._2954_ sky130_fd_sc_hd__nor2_1
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _05890_ _05889_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or2b_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3785_ MuI._2884_ vssd1 vssd1 vccd1 vccd1 MuI._2885_ sky130_fd_sc_hd__clkbuf_4
XMuI._6573_ MuI._2308_ MuI._2472_ vssd1 vssd1 vccd1 vccd1 MuI._2474_ sky130_fd_sc_hd__or2_1
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5113__D MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5524_ MuI._1313_ MuI._1317_ MuI._1319_ vssd1 vssd1 vccd1 vccd1 MuI._1320_ sky130_fd_sc_hd__nand3_1
X_07630_ _00228_ _00229_ _00246_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08541__A2 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._404_ AuI.pe.significand\[12\] AuI.pe.significand\[13\] AuI.pe.significand\[14\]
+ AuI.pe.significand\[15\] vssd1 vssd1 vccd1 vccd1 AuI.pe._371_ sky130_fd_sc_hd__or4_1
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5464__B2 MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5455_ MuI._1200_ MuI._1199_ MuI._1191_ vssd1 vssd1 vccd1 vccd1 MuI._1244_ sky130_fd_sc_hd__a21o_1
XFILLER_81_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5410__B MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1329_ AuI._0518_ AuI._0524_ vssd1 vssd1 vccd1 vccd1 AuI._0525_ sky130_fd_sc_hd__nand2_1
X_07561_ _00176_ _00177_ _00175_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__a21bo_1
XFILLER_207_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4406_ MuI._0087_ MuI._0089_ MuI.b_operand\[17\] MuI._3363_ vssd1 vssd1 vccd1
+ vccd1 MuI._0090_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ _02862_ _03906_ _01916_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5386_ MuI._1121_ MuI._1167_ vssd1 vssd1 vccd1 vccd1 MuI._1168_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07492_ net119 _00033_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__nand2_1
XFILLER_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4026__B MuI._0526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4337_ MuI._3387_ MuI._0009_ vssd1 vssd1 vccd1 vccd1 MuI._0015_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._1538__A AuI._0599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09231_ _01625_ _01674_ _01848_ _01437_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a211oi_2
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__A2_N _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10628__A _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__B1 _05126_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4268_ MuI._0614_ MuI._2830_ MuI._3247_ MuI._0361_ vssd1 vssd1 vccd1 vccd1 MuI._3368_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12546__C _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _01776_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__and2b_1
XANTENNA__09201__B _02194_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08743__D _00301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6007_ MuI._3094_ MuI._3096_ vssd1 vssd1 vccd1 vccd1 MuI._1851_ sky130_fd_sc_hd__nand2_1
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6241__B MuI._0537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ _00729_ _00730_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__nor2_1
XANTENNA__07002__A _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5519__A2 MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4199_ MuI._3291_ MuI._3290_ vssd1 vssd1 vccd1 vccd1 MuI._3299_ sky130_fd_sc_hd__or2b_1
XFILLER_147_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09093_ _01696_ _01708_ _01709_ _01710_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a211oi_4
XANTENNA__11600__A2 _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _00653_ _00656_ _00657_ _00658_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07937__A _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06841__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3950__A1 MuI._2055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09995_ _02660_ _02659_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__nand3_1
XANTENNA__13105__A2 _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__A2 _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _01547_ _01548_ _01562_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11116__A1 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07672__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13393__B _06016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _01492_ _01493_ _01494_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__nand3_2
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__A _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07391__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07828_ _00046_ _06605_ _06591_ _00049_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a22o_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5320__B MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4862__D MuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07759_ _00374_ _00375_ _00376_ vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__nand3_1
XFILLER_71_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10627__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08296__A1 _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _04133_ _02726_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__nor2_1
XFILLER_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12092__A2 _06546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _02048_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__and2b_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5758__A2 MuI._2341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _03539_ _03593_ _06518_ _00412_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__and4_1
XANTENNA__08048__A1 _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__A1 _02751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ _05201_ _05202_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__nor3b_4
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _03959_ _04054_ _04088_ _04089_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a211oi_4
XFILLER_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06751__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A1 _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _02760_ _03838_ _02192_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__o21a_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10273__A _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _02766_ _02880_ _02885_ _02761_ _02759_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a311o_1
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11184_ _03938_ _03940_ _03920_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._3941__D MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _03842_ _05992_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__and2_1
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08771__A2 _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11107__A1 _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10066_ _02738_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11658__A2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5511__A MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3570_ MuI._0966_ MuI._0933_ vssd1 vssd1 vccd1 vccd1 MuI._1626_ sky130_fd_sc_hd__or2b_1
XFILLER_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5230__B MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5240_ MuI._1003_ MuI._1006_ vssd1 vssd1 vccd1 vccd1 MuI._1007_ sky130_fd_sc_hd__xnor2_1
XAuI._1114_ AuI._0322_ AuI._0323_ vssd1 vssd1 vccd1 vccd1 AuI._0324_ sky130_fd_sc_hd__xor2_1
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10618__B1 _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06926__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ _03705_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__xnor2_4
XFILLER_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5171_ MuI._0885_ MuI._0893_ vssd1 vssd1 vccd1 vccd1 MuI._0931_ sky130_fd_sc_hd__or2b_1
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1045_ AuI._0256_ vssd1 vssd1 vccd1 vccd1 AuI._0257_ sky130_fd_sc_hd__buf_2
X_12707_ _05578_ _03186_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__B1 _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6342__A MuI._0372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._4122_ MuI._3219_ MuI._3221_ vssd1 vssd1 vccd1 vccd1 MuI._3222_ sky130_fd_sc_hd__or2b_1
X_10899_ _03460_ _03632_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__nand3b_2
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12638_ _00270_ _03449_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__nand2_1
XFILLER_129_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4421__A2 MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__B _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4053_ MuI._3125_ MuI._3152_ vssd1 vssd1 vccd1 vccd1 MuI._3153_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12085__D _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__A _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__xor2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07757__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07262__A2 _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07476__B _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4955_ MuI.b_operand\[10\] MuI._2837_ MuI.a_operand\[9\] MuI.a_operand\[8\] vssd1
+ vssd1 vccd1 vccd1 MuI._0694_ sky130_fd_sc_hd__and4_1
XFILLER_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4947__D MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0829_ AuI._0047_ AuI._0048_ vssd1 vssd1 vccd1 vccd1 AuI._0049_ sky130_fd_sc_hd__nor2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07195__C net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13494__A _06408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3906_ MuI._2996_ MuI._3004_ MuI._3005_ vssd1 vssd1 vccd1 vccd1 MuI._3006_ sky130_fd_sc_hd__and3_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _01416_ _01417_ _06608_ _00303_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__and4bb_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4886_ MuI._0616_ MuI._0617_ MuI._2796_ MuI._0101_ vssd1 vssd1 vccd1 vccd1 MuI._0618_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_140_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13099__A1 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _02426_ _02428_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__and2b_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _05338_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and3_1
XFILLER_140_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08588__A _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6625_ MuI._1413_ MuI._2530_ vssd1 vssd1 vccd1 vccd1 MuI._2531_ sky130_fd_sc_hd__xnor2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3837_ MuI._2935_ MuI._2936_ vssd1 vssd1 vccd1 vccd1 MuI._2937_ sky130_fd_sc_hd__xnor2_1
X_08731_ _06622_ _04574_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__nand2_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10630__B _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3768_ MuI.b_operand\[6\] vssd1 vssd1 vccd1 vccd1 MuI._2868_ sky130_fd_sc_hd__buf_2
XMuI._6556_ MuI._2452_ MuI._2454_ vssd1 vssd1 vccd1 vccd1 MuI._2455_ sky130_fd_sc_hd__and2_1
XANTENNA__08738__D _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08662_ _00975_ _00974_ _00973_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07642__D _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5507_ MuI._2967_ MuI._0315_ vssd1 vssd1 vccd1 vccd1 MuI._1301_ sky130_fd_sc_hd__nand2_1
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ net51 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__buf_2
XFILLER_81_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6487_ MuI._2377_ MuI._2371_ MuI._2376_ vssd1 vssd1 vccd1 vccd1 MuI._2379_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._5140__B MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3699_ MuI.b_operand\[13\] vssd1 vssd1 vccd1 vccd1 MuI._2799_ sky130_fd_sc_hd__buf_2
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _01204_ _01208_ _01210_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__o21a_1
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5438_ MuI._1223_ MuI._1224_ vssd1 vssd1 vccd1 vccd1 MuI._1225_ sky130_fd_sc_hd__nor2_1
X_07544_ _06480_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__buf_4
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06836__A _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3876__A MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5369_ MuI._1146_ MuI._1147_ MuI._1148_ vssd1 vssd1 vccd1 vccd1 MuI._1149_ sky130_fd_sc_hd__o21ba_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__A2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07475_ _04434_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__buf_6
XANTENNA_MuI._5794__C MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__inv_2
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09145_ _01753_ _01755_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__nor2_1
XFILLER_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _01685_ _01692_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08450__A1 _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08027_ _06576_ _06577_ _06639_ _06640_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__a22o_1
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10093__A _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08202__A1 _00162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08202__B2 _00164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _02634_ _02637_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__nor2_1
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4479__A2 MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08929_ _01495_ _01533_ _01545_ _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a211oi_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__B _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _04753_ _04754_ _04654_ _04602_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__o211a_2
XANTENNA__10848__B1 _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4592__D MuI._3246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _03324_ _05262_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__nand2_1
XFILLER_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _03363_ _03367_ _03548_ _03549_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__a211o_1
XFILLER_44_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10076__A1 _06428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3786__A MuI._2885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _03180_ _03279_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10268__A _00707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4939__B1 MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _02822_ _06367_ _02920_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ _03152_ _06605_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__and2_1
XFILLER_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09769__A1 _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _05272_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09769__B2 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6156__A2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ _05183_ _05107_ _05199_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a211oi_4
XFILLER_181_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11305_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__nor2_1
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _05124_ _05125_ _04987_ _04989_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a211o_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3914__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3914__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ _03822_ _03819_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__and2b_1
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1663_ AuI.exponent_sub\[5\] AuI._0599_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0016_
+ sky130_fd_sc_hd__o21a_1
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12930__B _05391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4740_ MuI.a_operand\[17\] MuI.a_operand\[16\] MuI.b_operand\[4\] MuI._2880_
+ vssd1 vssd1 vccd1 vccd1 MuI._0457_ sky130_fd_sc_hd__and4_1
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07645__A2_N _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11167_ _02754_ _02797_ _03424_ _00382_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and4_1
XAuI._1594_ AuI._0626_ AuI._0766_ vssd1 vssd1 vccd1 vccd1 AuI._0767_ sky130_fd_sc_hd__xor2_1
XFILLER_68_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4671_ MuI._1010_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0381_ sky130_fd_sc_hd__nand2_1
XFILLER_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _02862_ _04865_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__and2b_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11098_ _02751_ _03689_ _03835_ _03848_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__a211o_2
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__C _00359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__B _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6410_ MuI._2107_ MuI._2244_ MuI._2282_ vssd1 vssd1 vccd1 vccd1 MuI._2294_ sky130_fd_sc_hd__a21oi_1
XMuI._3622_ MuI._1780_ MuI._2165_ MuI._2132_ vssd1 vssd1 vccd1 vccd1 MuI._2198_ sky130_fd_sc_hd__or3b_1
XFILLER_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10049_ _02064_ _02706_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__or2_2
XFILLER_209_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07462__D _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6341_ MuI._0625_ MuI._1494_ MuI._2077_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._2218_
+ sky130_fd_sc_hd__a22oi_1
XMuI._3553_ MuI._0383_ MuI._0636_ MuI._0801_ MuI._1043_ vssd1 vssd1 vccd1 vccd1 MuI._1439_
+ sky130_fd_sc_hd__and4_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6092__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6092__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6272_ MuI._2140_ MuI._2141_ vssd1 vssd1 vccd1 vccd1 MuI._2142_ sky130_fd_sc_hd__xnor2_1
XFILLER_205_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3484_ MuI._0592_ MuI._0471_ MuI._0669_ MuI._0647_ vssd1 vssd1 vccd1 vccd1 MuI._0680_
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5223_ MuI._0986_ MuI._0987_ vssd1 vssd1 vccd1 vccd1 MuI._0989_ sky130_fd_sc_hd__or2_1
XFILLER_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3696__A MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10178__A _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__A2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0859__B2 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5154_ MuI._0873_ MuI._0875_ MuI._0874_ vssd1 vssd1 vccd1 vccd1 MuI._0913_ sky130_fd_sc_hd__o21bai_1
XAuI._1028_ net108 net124 net109 net125 AuI._0123_ AuI._0175_ vssd1 vssd1 vccd1 vccd1
+ AuI._0240_ sky130_fd_sc_hd__mux4_1
X_07260_ _06518_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__clkbuf_8
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4105_ MuI._3201_ MuI._3204_ vssd1 vssd1 vccd1 vccd1 MuI._3205_ sky130_fd_sc_hd__and2b_1
XANTENNA__08871__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5085_ MuI._0832_ MuI._0836_ vssd1 vssd1 vccd1 vccd1 MuI._0837_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._6222__D MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ _02096_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__buf_6
XFILLER_191_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5119__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08590__B _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4036_ MuI._1032_ MuI._1483_ MuI._2800_ MuI._2919_ vssd1 vssd1 vccd1 vccd1 MuI._3136_
+ sky130_fd_sc_hd__and4_1
XANTENNA__11567__B2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3862__C MuI._2874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _02532_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XMuI._5987_ MuI._1827_ MuI._1828_ vssd1 vssd1 vccd1 vccd1 MuI._1829_ sky130_fd_sc_hd__xnor2_1
XMuI._4938_ MuI._2440_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._0675_ sky130_fd_sc_hd__nand2_1
X_09832_ _02448_ _02482_ _02483_ _02443_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5658__A1 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._798_ AuI.pe._335_ AuI.pe._256_ AuI.pe._337_ AuI.pe._377_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._338_ sky130_fd_sc_hd__and4bb_1
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4869_ MuI._0597_ MuI._0595_ vssd1 vssd1 vccd1 vccd1 MuI._0599_ sky130_fd_sc_hd__xnor2_1
X_09763_ _00162_ _02409_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11456__B _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ _05155_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[18\] sky130_fd_sc_hd__clkbuf_2
XANTENNA__10360__B _06477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6608_ MuI._1795_ MuI._1808_ MuI._1831_ MuI._2511_ vssd1 vssd1 vccd1 vccd1 MuI._2512_
+ sky130_fd_sc_hd__a22oi_1
X_08714_ net110 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__buf_2
XFILLER_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08468__D _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _02333_ _02335_ _02330_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13492__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6539_ MuI._2405_ MuI._2435_ vssd1 vssd1 vccd1 vccd1 MuI._2436_ sky130_fd_sc_hd__nor2_1
XANTENNA__09160__A2 _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _01262_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08765__B _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13244__A1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _00941_ _00942_ _00943_ _00908_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__a22oi_2
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07527_ _00143_ _00142_ _06639_ _06637_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__o211a_1
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09299__D _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07458_ _00073_ _00075_ net114 _04240_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__and4bb_1
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3756__D MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07389_ _00004_ _00005_ _00006_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nand3_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12755__B1 _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09128_ _01743_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _01625_ _01622_ _01624_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__and3_1
XFILLER_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12507__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ _02844_ _04893_ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__o21a_1
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11021_ _00088_ _05036_ _03762_ _03763_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._4884__B MuI._2638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5061__A MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10701__D _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12972_ _05779_ _05828_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__nand2_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input11_A a_operand[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _04579_ _04583_ _04735_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a211oi_2
XANTENNA__09151__A2 _04638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0805__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A1 _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _06610_ _05777_ _04502_ _04501_ _05895_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__a32o_1
XFILLER_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4624__A2 MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0839__A_N net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__B2 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6604__B MuI._1836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10805_ _03530_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__nor2_2
XFILLER_202_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ _04460_ _04571_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__o211ai_2
XFILLER_198_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08111__B1 _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10736_ _03456_ _03457_ _03447_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a21o_1
XFILLER_202_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5585__B1 MuI._0111_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13455_ _02822_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__or2_1
X_10667_ _00444_ _05123_ _03382_ _03383_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a22o_1
XFILLER_51_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ AuI.result\[15\] _02938_ _05256_ _02935_ vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__D _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1266__A1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13386_ _06200_ _06201_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a31o_1
XFILLER_182_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ AuI.result\[2\] _02732_ _03308_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a211o_1
XMuI._5910_ MuI._1689_ MuI._1694_ vssd1 vssd1 vccd1 vccd1 MuI._1744_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._5236__A MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ _05071_ _05073_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or2b_1
XFILLER_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10772__A2 _02737_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5841_ MuI._1581_ MuI._1583_ MuI._1588_ vssd1 vssd1 vccd1 vccd1 MuI._1668_ sky130_fd_sc_hd__nor3b_1
XFILLER_5_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ _05105_ _05106_ _04965_ _04969_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o211ai_1
XAuI.pe._721_ AuI.pe._170_ AuI.pe._078_ AuI.pe._261_ AuI.pe._266_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._267_ sky130_fd_sc_hd__a211o_1
XMuI._5772_ MuI._1589_ MuI._1590_ MuI._1574_ vssd1 vssd1 vccd1 vccd1 MuI._1592_ sky130_fd_sc_hd__a21o_1
XFILLER_123_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _03966_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1646_ AuI.exp_a AuI.operand_a\[24\] AuI._0710_ AuI._0002_ vssd1 vssd1 vccd1
+ vccd1 AuI._0003_ sky130_fd_sc_hd__a31o_1
XFILLER_110_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12199_ _04951_ _04953_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__nor2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 ALU_Output[29] sky130_fd_sc_hd__buf_2
XAuI.pe._652_ AuI.pe._201_ AuI.pe._025_ AuI.pe._036_ vssd1 vssd1 vccd1 vccd1 AuI.pe._202_
+ sky130_fd_sc_hd__a21o_1
XMuI._4723_ MuI._0429_ MuI._0436_ MuI._0437_ vssd1 vssd1 vccd1 vccd1 MuI._0439_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._6301__A2 MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1577_ AuI._0259_ AuI._0751_ AuI._0752_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[10\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__C _00088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._583_ AuI.pe._056_ AuI.pe._086_ AuI.pe._137_ vssd1 vssd1 vccd1 vccd1 AuI.pe._138_
+ sky130_fd_sc_hd__a21o_1
XFILLER_95_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4654_ MuI._0360_ MuI._0362_ vssd1 vssd1 vccd1 vccd1 MuI._0363_ sky130_fd_sc_hd__nor2_1
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06760_ _02840_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__buf_8
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3605_ MuI._1989_ MuI._2000_ vssd1 vssd1 vccd1 vccd1 MuI._2011_ sky130_fd_sc_hd__and2b_1
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4585_ MuI._2803_ MuI._2786_ MuI._2352_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._0287_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_209_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06691_ _02096_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__buf_4
XFILLER_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5844__A2_N MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6324_ MuI._2157_ MuI._2140_ MuI._2141_ vssd1 vssd1 vccd1 vccd1 MuI._2200_ sky130_fd_sc_hd__or3b_1
XANTENNA__08585__B _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11292__A _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3536_ MuI._1230_ MuI._1241_ vssd1 vssd1 vccd1 vccd1 MuI._1252_ sky130_fd_sc_hd__and2_1
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12819__C _06537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ _01035_ _01046_ _01047_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__nand3_1
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6255_ MuI._2914_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._2124_ sky130_fd_sc_hd__nand2_1
XMuI._3467_ MuI.a_operand\[24\] MuI.a_operand\[23\] MuI.a_operand\[26\] MuI.a_operand\[25\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0493_ sky130_fd_sc_hd__nor4_4
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ _06504_ _05101_ _06517_ _06503_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__a22oi_1
XFILLER_211_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5206_ MuI._0967_ MuI._0968_ MuI._0965_ vssd1 vssd1 vccd1 vccd1 MuI._0970_ sky130_fd_sc_hd__a21o_1
X_07312_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__buf_6
XMuI._6186_ MuI._2813_ MuI._1483_ MuI._2066_ MuI._2814_ vssd1 vssd1 vccd1 vccd1 MuI._2048_
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08292_ _03454_ _03884_ _03982_ _03389_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12835__B _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5137_ MuI._0885_ MuI._0893_ vssd1 vssd1 vccd1 vccd1 MuI._0894_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ net108 vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__buf_4
XFILLER_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5068_ MuI._0816_ MuI._0817_ vssd1 vssd1 vccd1 vccd1 MuI._0818_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout129_A net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._3873__B MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ net108 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__clkbuf_8
XFILLER_180_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4019_ MuI._3103_ MuI._3104_ MuI._3118_ vssd1 vssd1 vccd1 vccd1 MuI._3119_ sky130_fd_sc_hd__or3_1
XANTENNA__07010__A _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6676__S MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4985__A MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12570__B _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input3_A Operation[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09815_ _02451_ _02452_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__and3_1
XFILLER_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _02387_ _02390_ _02391_ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a211oi_2
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06958_ _04972_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__buf_4
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11476__B1 _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _02187_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__xnor2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07144__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _04229_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08341__B1 _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07144__B2 _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08628_ _02754_ _02797_ _00083_ _00098_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__and4_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _01124_ _01131_ _01132_ _01176_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__o31a_1
XFILLER_196_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12976__B1 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _02604_ _02724_ _04351_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a211o_1
XFILLER_168_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ _06682_ _05509_ _05574_ _00000_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a22o_1
XFILLER_168_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ AuI.result\[25\] _02732_ _06145_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10452_ _03141_ _03142_ _03151_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5319__B1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ _02805_ _02809_ _05762_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or4_1
X_10383_ _03069_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__xor2_2
XFILLER_164_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ _04949_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__xnor2_2
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input59_A b_operand[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1500_ AuI._0678_ AuI._0681_ AuI._0684_ AuI._0685_ AuI._0679_ vssd1 vssd1 vccd1
+ vccd1 AuI._0686_ sky130_fd_sc_hd__o311ai_4
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ _04322_ _04874_ _04877_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__o21ba_1
XFILLER_132_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ _00058_ _06561_ _03743_ _03745_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__nand4_1
XAuI._1431_ AuI._0615_ AuI._0616_ vssd1 vssd1 vccd1 vccd1 AuI._0617_ sky130_fd_sc_hd__nand2_1
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07383__A1 _06682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__B2 _00000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1362_ AuI._0549_ AuI._0550_ vssd1 vssd1 vccd1 vccd1 AuI._0555_ sky130_fd_sc_hd__nand2_1
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _02805_ _05762_ _04211_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__o21a_1
XAuI._1293_ AuI._0486_ AuI._0490_ vssd1 vssd1 vccd1 vccd1 AuI._0492_ sky130_fd_sc_hd__nand2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4370_ MuI._0049_ MuI._0050_ vssd1 vssd1 vccd1 vccd1 MuI._0051_ sky130_fd_sc_hd__xnor2_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _04717_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nor2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _02751_ _05687_ _05688_ _05754_ _05771_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__a311o_4
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ MuI.result\[11\] _02738_ _04642_ _04607_ _04643_ vssd1 vssd1 vccd1 vccd1
+ _04644_ sky130_fd_sc_hd__a221o_1
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5270__A2 MuI._3402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6040_ MuI._0339_ MuI._2975_ vssd1 vssd1 vccd1 vccd1 MuI._1887_ sky130_fd_sc_hd__and2_2
XFILLER_199_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11768_ _04568_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__xnor2_4
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06934__A _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10719_ _03437_ _03438_ _03417_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__a21o_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08770__B_N _01387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _02860_ _04494_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__nand2_1
XFILLER_174_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13438_ _04161_ _06342_ _06343_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__a31o_1
XFILLER_127_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10175__B _05134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12093__D _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ _06279_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__nor2_1
XFILLER_170_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11942__A1 _04755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6873_ MuI._2772_ MuI._2498_ vssd1 vssd1 vccd1 vccd1 MuI._2774_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07765__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5824_ MuI._1573_ MuI._1631_ MuI._1632_ vssd1 vssd1 vccd1 vccd1 MuI._1650_ sky130_fd_sc_hd__nand3_1
XFILLER_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _00546_ _00547_ _06593_ _04843_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__and4bb_1
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._704_ AuI.pe._145_ AuI.pe._399_ AuI.pe._249_ AuI.pe._250_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._251_ sky130_fd_sc_hd__a211o_1
XFILLER_111_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5755_ MuI._1513_ MuI._1514_ MuI._1512_ vssd1 vssd1 vccd1 vccd1 MuI._1574_ sky130_fd_sc_hd__o21bai_1
XFILLER_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1629_ AuI._0681_ AuI._0794_ vssd1 vssd1 vccd1 vccd1 AuI._0795_ sky130_fd_sc_hd__xor2_1
X_07861_ _00438_ _00439_ _00477_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__and3_1
XFILLER_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._635_ AuI.pe._045_ AuI.pe._142_ AuI.pe._395_ vssd1 vssd1 vccd1 vccd1 AuI.pe._186_
+ sky130_fd_sc_hd__and3_1
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4706_ MuI._0321_ vssd1 vssd1 vccd1 vccd1 MuI._0420_ sky130_fd_sc_hd__clkbuf_4
X_09600_ _02170_ _02235_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__or2_1
XFILLER_56_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06812_ _03400_ _03121_ _03185_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__and3_1
XFILLER_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5686_ MuI._1490_ MuI._1491_ MuI._1497_ vssd1 vssd1 vccd1 vccd1 MuI._1498_ sky130_fd_sc_hd__nand3_1
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._5132__C MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07792_ _00173_ _00181_ _00180_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4836__A2 MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08596__A _01203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4029__B MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._566_ AuI.pe._028_ AuI.pe._112_ AuI.pe._119_ AuI.pe._030_ AuI.pe._121_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._122_ sky130_fd_sc_hd__a221o_1
XFILLER_49_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4637_ MuI.a_operand\[17\] MuI._2884_ MuI._3307_ MuI._1461_ vssd1 vssd1 vccd1
+ vccd1 MuI._0344_ sky130_fd_sc_hd__a22oi_1
X_09531_ _02138_ _02143_ _02159_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a211o_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06743_ _02658_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__buf_6
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._497_ AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 AuI.pe._059_ sky130_fd_sc_hd__clkbuf_4
XMuI._4568_ MuI._0104_ MuI._0098_ vssd1 vssd1 vccd1 vccd1 MuI._0268_ sky130_fd_sc_hd__and2b_1
X_09462_ _02052_ _02060_ _02073_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__and3_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07650__D _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6307_ MuI._2849_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._2181_ sky130_fd_sc_hd__nand2_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3519_ MuI._0383_ MuI._0636_ MuI._0592_ MuI._0801_ vssd1 vssd1 vccd1 vccd1 MuI._1065_
+ sky130_fd_sc_hd__and4_1
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08413_ _06630_ _04585_ _04649_ _06631_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__a22o_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4499_ MuI._0190_ MuI._0188_ vssd1 vssd1 vccd1 vccd1 MuI._0192_ sky130_fd_sc_hd__xnor2_1
X_09393_ _01907_ _01909_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11172__D _00785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6238_ MuI._0350_ MuI._2860_ MuI._2800_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._2105_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12958__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08344_ _00829_ _00828_ _00827_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06844__A _03744_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3884__A MuI._2843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6169_ MuI._0570_ MuI._2800_ MuI._2919_ MuI._0339_ vssd1 vssd1 vccd1 vccd1 MuI._2029_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08275_ _00890_ _00882_ _00889_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__and3_1
XFILLER_165_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07226_ _06519_ _06515_ net17 net18 vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__and4_1
XANTENNA__08481__D _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10085__B _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09874__B _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ _06452_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__and2_1
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0989__A0 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ _06356_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_161_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout110 net62 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_4
XFILLER_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout121 net42 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_6
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout132 net16 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13438__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ _02366_ _02372_ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nor3_2
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12459__C _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _05502_ _05505_ _05503_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o21bai_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._6154__B MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__A2 _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12671_ _05538_ _05539_ _05528_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5252__A2 MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _04409_ _04410_ _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__and3_1
XFILLER_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4460__B1 MuI.b_operand\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3794__A MuI._0559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09130__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ _02924_ _02775_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._6170__A MuI._0328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10707__C _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10504_ _03206_ _03207_ _03208_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and3_1
XFILLER_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0931_ AuI._0031_ AuI._0141_ AuI._0142_ AuI._0101_ vssd1 vssd1 vccd1 vccd1 AuI._0143_
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07288__C _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11484_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__and2_1
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12177__B2 _04736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ _06051_ _06050_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__and2_1
XFILLER_124_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _03831_ _04068_ _02975_ _02973_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__a31o_1
XFILLER_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0862_ net68 vssd1 vssd1 vccd1 vccd1 AuI._0082_ sky130_fd_sc_hd__inv_2
XFILLER_152_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _05908_ _05982_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__and2b_1
X_10366_ _03050_ _03059_ _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nand3_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10723__B _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _04931_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__and2b_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3870_ MuI._1032_ MuI._2898_ MuI._2902_ MuI._2900_ vssd1 vssd1 vccd1 vccd1 MuI._2970_
+ sky130_fd_sc_hd__a31o_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _05983_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ _00292_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__clkbuf_8
XFILLER_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12036_ _04813_ _04814_ _04856_ _04857_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__o22a_1
XFILLER_120_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5540_ MuI._2886_ MuI._2882_ MuI._0445_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._1337_
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11835__A _02944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1414_ AuI._0593_ AuI._0601_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[23\]
+ sky130_fd_sc_hd__xnor2_2
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._420_ AuI.pe.significand\[17\] AuI.pe._385_ AuI.pe._386_ AuI.pe.significand\[20\]
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._387_ sky130_fd_sc_hd__nor4_4
XANTENNA__06929__A _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5471_ MuI._2967_ MuI._0111_ MuI._1247_ MuI._1246_ vssd1 vssd1 vccd1 vccd1 MuI._1261_
+ sky130_fd_sc_hd__a31o_1
XFILLER_207_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1345_ AuI._0524_ AuI._0537_ vssd1 vssd1 vccd1 vccd1 AuI._0540_ sky130_fd_sc_hd__nor2_1
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4422_ MuI.b_operand\[22\] MuI.b_operand\[21\] MuI._3247_ MuI._3372_ vssd1 vssd1
+ vccd1 vccd1 MuI._0107_ sky130_fd_sc_hd__and4_1
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1276_ AuI._0466_ AuI._0473_ AuI._0475_ vssd1 vssd1 vccd1 vccd1 AuI._0476_ sky130_fd_sc_hd__a21oi_4
X_12938_ _05780_ _05781_ _05825_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__or3_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4353_ MuI._0028_ MuI._0031_ vssd1 vssd1 vccd1 vccd1 MuI._0033_ sky130_fd_sc_hd__xnor2_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _05748_ _05752_ _06428_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a21oi_1
XMuI._4284_ MuI._3340_ MuI._3380_ MuI._3381_ vssd1 vssd1 vccd1 vccd1 MuI._3384_ sky130_fd_sc_hd__or3b_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6023_ MuI._1864_ MuI._1867_ vssd1 vssd1 vccd1 vccd1 MuI._1869_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07479__B _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6080__A MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ net57 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_2
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07011_ _05542_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[24\] sky130_fd_sc_hd__clkbuf_2
XFILLER_174_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11729__B _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5424__A MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6856_ MuI.b_operand\[23\] MuI._2489_ vssd1 vssd1 vccd1 vccd1 MuI._2760_ sky130_fd_sc_hd__xnor2_1
X_08962_ _01208_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__nor2_1
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5807_ MuI._1541_ MuI._1543_ MuI._1629_ MuI._1630_ vssd1 vssd1 vccd1 vccd1 MuI._1631_
+ sky130_fd_sc_hd__a211o_1
X_07913_ _00162_ _00412_ _00530_ _00164_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__a22oi_2
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6787_ MuI._2563_ MuI._2509_ MuI._2486_ vssd1 vssd1 vccd1 vccd1 MuI._2709_ sky130_fd_sc_hd__mux2_1
XMuI._3999_ MuI._3096_ MuI._3097_ MuI._3092_ vssd1 vssd1 vccd1 vccd1 MuI._3099_ sky130_fd_sc_hd__a21o_1
X_08893_ _01358_ _01363_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__and2_1
XANTENNA__11167__D _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12340__A1 _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1396__A0 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5738_ MuI._1464_ MuI._1554_ vssd1 vssd1 vccd1 vccd1 MuI._1555_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07844_ net117 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__buf_4
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06839__A _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._618_ AuI.pe.significand\[14\] vssd1 vssd1 vccd1 vccd1 AuI.pe._170_ sky130_fd_sc_hd__buf_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08757__C _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5669_ MuI._1014_ MuI._1015_ MuI._1052_ MuI._1053_ vssd1 vssd1 vccd1 vccd1 MuI._1479_
+ sky130_fd_sc_hd__nor4_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07775_ _00389_ _00391_ _00390_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__a21o_1
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6255__A MuI._2914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._549_ AuI.pe._105_ vssd1 vssd1 vccd1 vccd1 AuI.pe._106_ sky130_fd_sc_hd__buf_2
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ _02087_ _02139_ _02141_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__or4_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06726_ _02474_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__buf_4
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09445_ _02062_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09376_ _01939_ _01941_ _01942_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__and3_1
XFuI._100_ FuI._052_ FuI._059_ FuI.a_operand\[9\] vssd1 vssd1 vccd1 vccd1 FuI._021_
+ sky130_fd_sc_hd__o21a_1
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12295__B _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08327_ _00653_ _00654_ _00620_ _00655_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a22oi_2
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08075__A2 _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08258_ _00011_ _00048_ _00040_ _00012_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__a22o_1
XANTENNA_MuI._5318__B MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07209_ _06473_ _06474_ _06484_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21o_1
XFILLER_193_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08189_ _00712_ _00806_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__xnor2_2
XFILLER_180_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _02901_ _02856_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a21o_1
XANTENNA__12742__C _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _02827_ _05724_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__and2_1
XFILLER_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5053__B MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _02715_ _02753_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07889__A2 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06749__A _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09770__D net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1130_ AuI._0206_ AuI._0236_ AuI._0279_ AuI._0338_ vssd1 vssd1 vccd1 vccd1 AuI._0339_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._3484__A1 MuI._0592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ _03721_ _03723_ _03724_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__a21o_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10645__A1 _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ _02868_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__nand2_1
XAuI._1061_ AuI._0164_ AuI._0169_ AuI._0218_ vssd1 vssd1 vccd1 vccd1 AuI._0272_ sky130_fd_sc_hd__and3_1
XFILLER_204_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07510__A1 _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12917__C _05585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ _05429_ _05430_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__and2_1
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3787__A2 MuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11605_ _04392_ _04393_ _04394_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__a21o_1
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07299__B _06599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__D _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12585_ _00283_ _06546_ _05447_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__a22o_1
XFILLER_184_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._6186__B1 MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ _03664_ _04314_ _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a21o_1
XFILLER_157_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._0914_ AuI._0132_ vssd1 vssd1 vccd1 vccd1 AuI.operand_a\[24\] sky130_fd_sc_hd__clkbuf_2
XFILLER_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _04244_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__or2_1
XFILLER_109_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _02815_ _06017_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nor2_1
XMuI._4971_ MuI._2918_ MuI._2319_ MuI._2829_ MuI._2799_ vssd1 vssd1 vccd1 vccd1 MuI._0711_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_171_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ _03113_ _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__xnor2_1
XFILLER_171_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11549__B _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0845_ net110 AuI._0062_ AuI._0047_ AuI._0048_ AuI._0064_ vssd1 vssd1 vccd1 vccd1
+ AuI._0065_ sky130_fd_sc_hd__a2111o_1
X_11398_ _04161_ _04164_ _04171_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__a21o_1
XMuI._6710_ MuI._2364_ MuI._2623_ vssd1 vssd1 vccd1 vccd1 MuI._2624_ sky130_fd_sc_hd__or2b_1
XFILLER_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3922_ MuI._2787_ MuI._2407_ MuI._3021_ vssd1 vssd1 vccd1 vccd1 MuI._3022_ sky130_fd_sc_hd__a21bo_1
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ _06036_ _06038_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _03005_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__xor2_2
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6641_ MuI._2547_ MuI._1236_ vssd1 vssd1 vccd1 vccd1 MuI._2548_ sky130_fd_sc_hd__nor2_1
XFILLER_140_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3853_ MuI._2926_ MuI._2952_ vssd1 vssd1 vccd1 vccd1 MuI._2953_ sky130_fd_sc_hd__xor2_1
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _05964_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nand2_1
XFILLER_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6572_ MuI._1758_ MuI._2297_ vssd1 vssd1 vccd1 vccd1 MuI._2472_ sky130_fd_sc_hd__and2_1
X_12019_ _04837_ _04838_ _04834_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a21o_1
XMuI._3784_ MuI.b_operand\[4\] vssd1 vssd1 vccd1 vccd1 MuI._2884_ sky130_fd_sc_hd__buf_2
XFILLER_93_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5523_ MuI._1295_ MuI._1297_ MuI._1312_ vssd1 vssd1 vccd1 vccd1 MuI._1319_ sky130_fd_sc_hd__a21o_1
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09035__A _01203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._403_ AuI.pe._367_ AuI.pe._368_ AuI.pe._369_ vssd1 vssd1 vccd1 vccd1 AuI.pe._370_
+ sky130_fd_sc_hd__or3_4
XFILLER_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5464__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5454_ MuI._1200_ MuI._1191_ MuI._1199_ vssd1 vssd1 vccd1 vccd1 MuI._1243_ sky130_fd_sc_hd__nand3_1
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1328_ AuI._0523_ vssd1 vssd1 vccd1 vccd1 AuI._0524_ sky130_fd_sc_hd__inv_2
X_07560_ _00175_ _00176_ _00177_ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__nand3b_1
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4405_ MuI._1791_ MuI._3349_ MuI._0088_ MuI._3000_ vssd1 vssd1 vccd1 vccd1 MuI._0089_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5385_ MuI._1157_ MuI._1166_ vssd1 vssd1 vccd1 vccd1 MuI._1167_ sky130_fd_sc_hd__nor2_1
X_07491_ net120 net44 _06611_ _06602_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__and4_1
XAuI._1259_ AuI._0457_ AuI._0459_ AuI._0455_ vssd1 vssd1 vccd1 vccd1 AuI._0460_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4336_ MuI._3304_ MuI._0013_ vssd1 vssd1 vccd1 vccd1 MuI._0014_ sky130_fd_sc_hd__nand2_1
X_09230_ _01626_ _01672_ _01673_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__nor3_2
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10628__B _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4267_ MuI._3360_ MuI._3366_ vssd1 vssd1 vccd1 vccd1 MuI._3367_ sky130_fd_sc_hd__xnor2_1
X_09161_ _01776_ _01777_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__or3_1
XANTENNA__13004__B _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6006_ MuI._3142_ MuI._3145_ vssd1 vssd1 vccd1 vccd1 MuI._1850_ sky130_fd_sc_hd__nand2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10939__A2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _03228_ _03282_ _04585_ _04649_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__and4_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4198_ MuI._3296_ MuI._3297_ vssd1 vssd1 vccd1 vccd1 MuI._3298_ sky130_fd_sc_hd__nand2_1
X_09092_ _01605_ _01606_ _01607_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__and3_1
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ _00588_ _00621_ _00659_ _00660_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__o211a_1
XFILLER_163_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07937__B _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout111_A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10644__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08114__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3950__A2 MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09994_ _02657_ _02656_ _02655_ _02650_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a211o_1
XFILLER_89_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6839_ MuI._2692_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2752_ sky130_fd_sc_hd__and2b_1
XANTENNA__07953__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08945_ _01560_ _01561_ _01549_ _01550_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a211o_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1369__B1 AuI._0560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08876_ _01485_ _01486_ _01491_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a21o_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _06603_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__buf_6
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07758_ _02205_ _00153_ net29 _06534_ vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__a22o_1
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5320__C MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__A _01394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06709_ _02291_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__buf_4
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10627__A1 _03615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _00284_ _00306_ vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__nor2_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08296__A2 _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _06515_ net124 net123 _06519_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _01971_ _01972_ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a21o_1
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08048__A2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__xnor2_2
XFILLER_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _04086_ _04087_ _03938_ _03941_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__o211a_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11252_ _04327_ _02727_ _02945_ _04262_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09548__A2 _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10273__B _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10203_ _02767_ _02882_ _02883_ _02884_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a211o_1
XFILLER_122_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _03920_ _03938_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand3_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10134_ _02783_ _02791_ _02810_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__or3b_1
XANTENNA_input41_A b_operand[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11107__A2 _04327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10065_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5511__B MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07731__A1 _03486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1113_ net27 net59 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0323_ sky130_fd_sc_hd__mux2_1
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _03706_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__clkinv_2
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10729__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5170_ MuI._0886_ MuI._0892_ vssd1 vssd1 vccd1 vccd1 MuI._0930_ sky130_fd_sc_hd__or2b_1
XFILLER_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _03024_ _05058_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__nor2_1
XAuI._1044_ AuI._0255_ vssd1 vssd1 vccd1 vccd1 AuI._0256_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11291__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _02388_ _05970_ _03630_ _03631_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__a22o_1
XMuI._4121_ MuI._3220_ MuI._2793_ vssd1 vssd1 vccd1 vccd1 MuI._3221_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._6342__B MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08791__A1_N _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12637_ _05502_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XFILLER_169_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4052_ MuI._3149_ MuI._3151_ vssd1 vssd1 vccd1 vccd1 MuI._3152_ sky130_fd_sc_hd__xor2_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12240__B1 _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ _03525_ _05198_ _05294_ _05293_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__a31o_1
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06942__A _04800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__B _05520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _04142_ _04145_ _04300_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__o211a_2
XANTENNA__07757__B net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._145__151 vssd1 vssd1 vccd1 vccd1 FuI._145__151/HI net151 sky130_fd_sc_hd__conb_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12499_ _04873_ _05352_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10183__B _02970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4954_ MuI._0682_ MuI._0689_ MuI._0692_ vssd1 vssd1 vccd1 vccd1 MuI._0693_ sky130_fd_sc_hd__a21o_1
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0828_ net124 net108 vssd1 vssd1 vccd1 vccd1 AuI._0048_ sky130_fd_sc_hd__and2b_1
XFILLER_140_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07195__D _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3905_ MuI._3002_ MuI._3003_ MuI._2997_ vssd1 vssd1 vccd1 vccd1 MuI._3005_ sky130_fd_sc_hd__a21o_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4885_ MuI._2803_ MuI._2374_ MuI._3363_ MuI._2802_ vssd1 vssd1 vccd1 vccd1 MuI._0617_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _05327_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__13099__A2 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6624_ MuI._1436_ MuI._1443_ MuI._1426_ vssd1 vssd1 vccd1 vccd1 MuI._2530_ sky130_fd_sc_hd__a21oi_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3836_ MuI._2748_ MuI._2783_ vssd1 vssd1 vccd1 vccd1 MuI._2936_ sky130_fd_sc_hd__and2_1
XFILLER_112_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08730_ _02712_ _04445_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__nand2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__B _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6555_ MuI._2449_ MuI._2453_ vssd1 vssd1 vccd1 vccd1 MuI._2454_ sky130_fd_sc_hd__nor2_1
XFILLER_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3767_ MuI._2866_ vssd1 vssd1 vccd1 vccd1 MuI._2867_ sky130_fd_sc_hd__clkbuf_4
X_08661_ _00975_ _00973_ _00974_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__or3_1
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5506_ MuI._1298_ MuI._1299_ vssd1 vssd1 vccd1 vccd1 MuI._1300_ sky130_fd_sc_hd__nor2_1
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07612_ net50 net51 _04509_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__and3_1
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6486_ MuI._2371_ MuI._2376_ MuI._2377_ vssd1 vssd1 vccd1 vccd1 MuI._2378_ sky130_fd_sc_hd__a21oi_2
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3698_ MuI._2796_ MuI._2797_ vssd1 vssd1 vccd1 vccd1 MuI._2798_ sky130_fd_sc_hd__nand2_1
X_08592_ _01160_ _01209_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__nor2_2
XANTENNA__08744__A1_N _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5437_ MuI._1218_ MuI._1220_ MuI._1222_ vssd1 vssd1 vccd1 vccd1 MuI._1224_ sky130_fd_sc_hd__and3_1
XFILLER_207_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07543_ _02291_ _06548_ _05627_ net130 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__and4_1
XFILLER_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10639__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5368_ MuI._2867_ MuI._2869_ MuI._3371_ MuI._0444_ vssd1 vssd1 vccd1 vccd1 MuI._1148_
+ sky130_fd_sc_hd__and4_1
XFILLER_210_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07474_ _00080_ _00091_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__nor2_1
XFILLER_195_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08109__A _00231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4319_ MuI._3277_ MuI._3276_ vssd1 vssd1 vccd1 vccd1 MuI._3419_ sky130_fd_sc_hd__and2b_1
XFILLER_167_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ _01825_ _01828_ _01829_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07013__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5299_ MuI._0810_ MuI._1071_ vssd1 vssd1 vccd1 vccd1 MuI._1072_ sky130_fd_sc_hd__and2b_1
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ _01735_ _01758_ _01760_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07948__A _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06852__A _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0900__B net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ _01686_ _01691_ _01687_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nand3_1
XFILLER_190_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08450__A2 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__B1 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08026_ _00641_ _00642_ _00561_ _00643_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__and4bb_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__B _04057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12534__A1 _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08202__A2 _06518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__A net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07683__A _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09977_ _02639_ _02641_ _01847_ _01881_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o211a_1
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08928_ _01537_ _01538_ _01544_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__and3_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__C _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10848__A1 _00096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10848__B2 _00095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__and2b_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4228__A MuI._2616_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _04677_ _04678_ _04679_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o21a_1
XANTENNA_MuI._5050__C MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _03546_ _03547_ _03536_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10549__A _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _03278_ _03276_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__and2b_1
XFILLER_125_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10268__B _00708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4939__A1 MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5059__A MuI._2873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4939__B2 MuI._2605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ _02814_ _02820_ _06365_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__or3_1
XFILLER_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10683_ _00133_ _00132_ _06591_ _06584_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__nand4_1
XFILLER_186_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12422_ _00270_ _03071_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__nand2_1
XANTENNA__09769__A2 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._129__135 vssd1 vssd1 vccd1 vccd1 FuI._129__135/HI net135 sky130_fd_sc_hd__conb_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06762__A _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_AuI._0810__B net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6220__A2_N MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__B1 _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12353_ _05196_ _05197_ _05099_ _05104_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__o211a_1
XFILLER_166_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ _03228_ _03282_ _05036_ _00534_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__and4_1
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12284_ _04987_ _04989_ _05124_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__o211ai_4
XANTENNA_AuI.pe._757__B2 AuI.pe.significand\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ _03861_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__xnor2_4
XAuI._1662_ AuI._0604_ AuI._0692_ AuI.operand_a\[28\] AuI._0258_ vssd1 vssd1 vccd1
+ vccd1 AuI._0015_ sky130_fd_sc_hd__a211o_1
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._509__A1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ _00878_ _05574_ _05649_ _00877_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a22oi_1
XAuI._1593_ AuI._0623_ AuI._0624_ AuI._0755_ AuI._0627_ vssd1 vssd1 vccd1 vccd1 AuI._0766_
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4670_ MuI._0376_ MuI._0379_ vssd1 vssd1 vccd1 vccd1 MuI._0380_ sky130_fd_sc_hd__nor2_1
XFILLER_67_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10117_ _04865_ _02862_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__and2b_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11097_ _02552_ _03315_ _03837_ _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a31o_1
XFILLER_110_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12004__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3621_ MuI._1494_ MuI._0471_ MuI._1450_ MuI._1439_ vssd1 vssd1 vccd1 vccd1 MuI._2187_
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10048_ _02718_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__buf_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6340_ MuI._2215_ MuI._2216_ vssd1 vssd1 vccd1 vccd1 MuI._2217_ sky130_fd_sc_hd__xnor2_1
XMuI._3552_ MuI._0636_ MuI._0801_ MuI._1043_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._1428_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6271_ MuI._2043_ MuI._2063_ vssd1 vssd1 vccd1 vccd1 MuI._2141_ sky130_fd_sc_hd__or2b_1
XANTENNA__09313__A net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3483_ MuI._0647_ MuI._0658_ vssd1 vssd1 vccd1 vccd1 MuI._0669_ sky130_fd_sc_hd__nor2_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5222_ MuI._1813_ MuI._0421_ MuI._0985_ vssd1 vssd1 vccd1 vccd1 MuI._0987_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _00421_ _04817_ _04818_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a21bo_1
XFILLER_189_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5153_ MuI._0909_ MuI._0910_ vssd1 vssd1 vccd1 vccd1 MuI._0912_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1027_ AuI._0237_ AuI._0238_ AuI._0031_ vssd1 vssd1 vccd1 vccd1 AuI._0239_ sky130_fd_sc_hd__mux2_1
XFILLER_177_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4104_ MuI._3202_ MuI._3203_ vssd1 vssd1 vccd1 vccd1 MuI._3204_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08871__B _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5084_ MuI._0833_ MuI._0835_ vssd1 vssd1 vccd1 vccd1 MuI._0836_ sky130_fd_sc_hd__xnor2_1
X_07190_ net116 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__buf_6
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4035_ MuI._2077_ MuI._2583_ vssd1 vssd1 vccd1 vccd1 MuI._3135_ sky130_fd_sc_hd__nand2_1
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5119__D MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07640__B1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3862__D MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _02118_ _03895_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__nand2_2
XMuI._5986_ MuI._1818_ MuI._1822_ vssd1 vssd1 vccd1 vccd1 MuI._1828_ sky130_fd_sc_hd__xnor2_1
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10922__A _03509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4937_ MuI.a_operand\[15\] MuI.a_operand\[14\] MuI._2884_ MuI._2880_ vssd1 vssd1
+ vccd1 vccd1 MuI._0674_ sky130_fd_sc_hd__and4_1
XFILLER_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09831_ _02448_ _02482_ _02483_ _02443_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__or4bb_1
XFILLER_112_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5658__A2 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._797_ AuI.pe._149_ AuI.pe._367_ AuI.pe._336_ AuI.pe._372_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._337_ sky130_fd_sc_hd__or4_1
XFILLER_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4868_ MuI._0595_ MuI._0597_ vssd1 vssd1 vccd1 vccd1 MuI._0598_ sky130_fd_sc_hd__and2b_1
XFILLER_101_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06974_ _05134_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__and3_1
X_09762_ _06480_ net127 net126 _06479_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a22o_1
XMuI._6607_ MuI._2510_ vssd1 vssd1 vccd1 vccd1 MuI._2511_ sky130_fd_sc_hd__inv_2
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3819_ MuI._2918_ vssd1 vssd1 vccd1 vccd1 MuI._2919_ sky130_fd_sc_hd__clkbuf_4
X_08713_ _00955_ _00956_ _01322_ _01327_ _01330_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o2111a_1
XANTENNA__07008__A _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4799_ MuI._0395_ MuI._0392_ MuI._0393_ vssd1 vssd1 vccd1 vccd1 MuI._0522_ sky130_fd_sc_hd__a21oi_1
X_09693_ _02330_ _02333_ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__and3_2
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6538_ MuI._2401_ MuI._2402_ MuI._2404_ vssd1 vssd1 vccd1 vccd1 MuI._2435_ sky130_fd_sc_hd__nor3_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _01252_ _01258_ _01261_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__a21oi_2
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6469_ MuI._2353_ MuI._2357_ MuI._2358_ vssd1 vssd1 vccd1 vccd1 MuI._2359_ sky130_fd_sc_hd__o21ba_1
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MuI._4094__A1 MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _01175_ _01177_ _01178_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__or3_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _06637_ _06639_ _00142_ _00143_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a211oi_4
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__B2 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10088__B _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__A1 _00734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _03271_ _00074_ _04358_ _03217_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12584__A _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0911__A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _02723_ _05047_ _06625_ _06624_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a31o_1
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ _01740_ _01742_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__nand2_1
XANTENNA__12755__A1 _00676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__B2 _00506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ _01437_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__xnor2_2
XANTENNA__10230__A2 _05724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08009_ _02107_ _06495_ _05434_ _06466_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__and4_1
XFILLER_117_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10832__A _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__A1 _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _00262_ _00421_ _03762_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nand4_1
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08302__A _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__B1 _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4884__C MuI._0088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A1_N _06439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5061__B MuI._3371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _02908_ _05860_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
XFILLER_58_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__B1_N _03186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _04733_ _04734_ _04723_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11494__A1 _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06757__A _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ _04659_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A2 _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12176__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10804_ _03517_ _03519_ _03529_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__and3_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _04584_ _04586_ _04454_ _04459_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__o211ai_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08111__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08111__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10735_ _03447_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__nand3_1
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4124__C MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5585__A1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ _06367_ _06368_ _02926_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__mux2_1
X_10666_ _00217_ _00216_ _00002_ _06568_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__nand4_1
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _05249_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__xnor2_1
X_13385_ _06200_ _06201_ _06270_ _06271_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a311o_1
X_10597_ _04133_ _02718_ _02721_ _02259_ _03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a221o_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5236__B MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _05092_ _05110_ _05109_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a21boi_2
XFILLER_182_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5840_ MuI._1665_ MuI._1666_ vssd1 vssd1 vccd1 vccd1 MuI._1667_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _04965_ _04969_ _05105_ _05106_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__a211o_2
XAuI.pe._720_ AuI.pe._142_ AuI.pe._112_ AuI.pe._264_ AuI.pe._265_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._266_ sky130_fd_sc_hd__a211o_1
XFILLER_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5771_ MuI._1574_ MuI._1589_ MuI._1590_ vssd1 vssd1 vccd1 vccd1 MuI._1591_ sky130_fd_sc_hd__nand3_1
X_11218_ _03976_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__or2b_1
XANTENNA_output72_A net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1645_ AuI.exponent_sub\[1\] AuI._0769_ AuI._0699_ vssd1 vssd1 vccd1 vccd1 AuI._0002_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_123_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12198_ _05024_ _05027_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__nor3_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._651_ AuI.pe._367_ vssd1 vssd1 vccd1 vccd1 AuI.pe._201_ sky130_fd_sc_hd__buf_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 ALU_Output[1] sky130_fd_sc_hd__buf_2
XMuI._4722_ MuI._0296_ MuI._0298_ vssd1 vssd1 vccd1 vccd1 MuI._0437_ sky130_fd_sc_hd__xnor2_1
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 ALU_Output[2] sky130_fd_sc_hd__buf_2
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11149_ _03900_ _03901_ _03774_ _03776_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__a211o_1
XAuI._1576_ AuI.pe.Significand\[10\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0752_
+ sky130_fd_sc_hd__or2_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07473__D _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._582_ AuI.pe._071_ AuI.pe._066_ AuI.pe._054_ AuI.pe._089_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._137_ sky130_fd_sc_hd__a22o_1
XFILLER_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4653_ MuI._0349_ MuI._0357_ MuI._0359_ vssd1 vssd1 vccd1 vccd1 MuI._0362_ sky130_fd_sc_hd__and3_1
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3604_ MuI._1978_ MuI._1923_ MuI._1956_ vssd1 vssd1 vccd1 vccd1 MuI._2000_ sky130_fd_sc_hd__or3_1
XANTENNA__11573__A _04302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4584_ MuI._2796_ MuI._2374_ vssd1 vssd1 vccd1 vccd1 MuI._0286_ sky130_fd_sc_hd__nand2_1
X_06690_ net37 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__buf_4
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6323_ MuI._2195_ MuI._2197_ vssd1 vssd1 vccd1 vccd1 MuI._2199_ sky130_fd_sc_hd__or2b_1
XFILLER_52_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3535_ MuI._1131_ MuI._1219_ vssd1 vssd1 vccd1 vccd1 MuI._1241_ sky130_fd_sc_hd__or2_1
XANTENNA__08585__C _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__B _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12819__D _05756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6254_ MuI._2849_ MuI._2120_ MuI._2122_ vssd1 vssd1 vccd1 vccd1 MuI._2123_ sky130_fd_sc_hd__a21bo_1
XFILLER_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3466_ MuI.a_operand\[28\] MuI.a_operand\[27\] MuI.a_operand\[29\] MuI.a_operand\[30\]
+ vssd1 vssd1 vccd1 vccd1 MuI._0482_ sky130_fd_sc_hd__nor4_4
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ net108 _05025_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__nand2_1
XMuI._5205_ MuI._0965_ MuI._0967_ MuI._0968_ vssd1 vssd1 vccd1 vccd1 MuI._0969_ sky130_fd_sc_hd__nand3_1
XFILLER_189_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07311_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__buf_4
XMuI._6185_ MuI._2939_ MuI._1142_ MuI._1483_ MuI._2066_ vssd1 vssd1 vccd1 vccd1 MuI._2047_
+ sky130_fd_sc_hd__and4_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08291_ _00610_ _00611_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5136_ MuI._0886_ MuI._0892_ vssd1 vssd1 vccd1 vccd1 MuI._0893_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07242_ _06539_ _06541_ _06540_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__a21o_1
XANTENNA__12835__C _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5067_ MuI._2838_ MuI._3245_ MuI._0304_ MuI._2836_ vssd1 vssd1 vccd1 vccd1 MuI._0817_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07173_ _06465_ _06472_ _06471_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a21o_1
XFILLER_192_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4018_ MuI._3111_ MuI._3117_ vssd1 vssd1 vccd1 vccd1 MuI._3118_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4985__B MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5969_ MuI._1795_ MuI._1808_ vssd1 vssd1 vccd1 vccd1 MuI._1809_ sky130_fd_sc_hd__xor2_1
XFILLER_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6258__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09814_ _02458_ _02464_ _02465_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a21o_1
XFILLER_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09745_ _02315_ _02314_ _02287_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a21oi_1
X_06957_ _04961_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__buf_4
XFILLER_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _02217_ _02215_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__and2b_1
X_06888_ net124 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__clkbuf_4
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__A2 _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _01228_ _01242_ _01243_ _01244_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__a211oi_4
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__A _01407_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08558_ _01120_ _01065_ _01122_ _00871_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__a211o_1
XFILLER_52_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__A1 _03454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__B2 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ _00125_ _00090_ _04445_ _00124_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__a22o_1
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ _01075_ _01076_ _01070_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__a21bo_1
XFILLER_195_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10827__A _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10520_ _03222_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__xnor2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _03149_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__xor2_1
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5319__A1 MuI._3349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13170_ _02779_ _02782_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__or2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10382_ _03076_ _03077_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__and2b_1
XFILLER_191_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ net60 _04918_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__and2_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4542__A2 MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _04614_ _04616_ _04761_ _04875_ _04760_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__o311ai_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__B _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6168__A MuI._0790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _03002_ _06561_ _03743_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a22o_1
XAuI._1430_ AuI._0560_ AuI._0557_ vssd1 vssd1 vccd1 vccd1 AuI._0616_ sky130_fd_sc_hd__or2b_1
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07383__A2 _06525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1361_ AuI._0551_ AuI._0554_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[18\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_93_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0816__A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _05843_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_2
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1292_ AuI._0486_ AuI._0490_ vssd1 vssd1 vccd1 vccd1 AuI._0491_ sky130_fd_sc_hd__or2_1
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11905_ _04705_ _04706_ _04716_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__and3_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05757_ _05758_ _05764_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a211o_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _04671_ _02941_ _02871_ _03306_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__o22ai_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12967__A1 _02801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _00502_ _04660_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__nand2_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10718_ _03417_ _03437_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand3_2
XFILLER_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11698_ _02860_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or2_1
XANTENNA__12719__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _03314_ _06345_ _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a21o_1
X_10649_ _03161_ _03164_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__nand2_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06950__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ _06231_ _06234_ _06278_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor3_1
XFILLER_182_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6872_ MuI._2499_ MuI._0207_ vssd1 vssd1 vccd1 vccd1 MuI._2772_ sky130_fd_sc_hd__and2b_1
XANTENNA__11942__A2 _04756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__B _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__xnor2_1
X_13299_ _02743_ _02831_ _02944_ _05595_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a22o_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4344__A_N MuI._0019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5823_ MuI._1473_ MuI._1572_ MuI._1569_ vssd1 vssd1 vccd1 vccd1 MuI._1649_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09348__B1 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._703_ AuI.pe._170_ AuI.pe._002_ AuI.pe._053_ AuI.pe._120_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._250_ sky130_fd_sc_hd__a22o_1
XFILLER_123_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5754_ MuI._1473_ MuI._1572_ vssd1 vssd1 vccd1 vccd1 MuI._1573_ sky130_fd_sc_hd__xor2_1
XAuI._1628_ AuI._0678_ AuI._0684_ AuI._0682_ vssd1 vssd1 vccd1 vccd1 AuI._0794_ sky130_fd_sc_hd__o21ba_1
X_07860_ _00438_ _00439_ _00477_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._634_ AuI.pe._120_ AuI.pe._184_ AuI.pe._141_ AuI.pe._372_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._185_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4705_ MuI._0375_ MuI._0414_ vssd1 vssd1 vccd1 vccd1 MuI._0419_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07781__A _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5685_ MuI._1495_ MuI._1496_ vssd1 vssd1 vccd1 vccd1 MuI._1497_ sky130_fd_sc_hd__xor2_1
XFILLER_56_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06811_ _03389_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__buf_4
XAuI._1559_ AuI._0736_ AuI._0737_ vssd1 vssd1 vccd1 vccd1 AuI._0738_ sky130_fd_sc_hd__nor2_1
X_07791_ _00407_ _00406_ _00185_ _00373_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a211o_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._565_ AuI.pe._033_ AuI.pe._120_ AuI.pe._388_ vssd1 vssd1 vccd1 vccd1 AuI.pe._121_
+ sky130_fd_sc_hd__and3_1
XANTENNA__08596__B _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09103__A2_N _04122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4636_ MuI._2840_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._0343_ sky130_fd_sc_hd__nand2_1
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4029__C MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _02147_ _02148_ _02157_ _02158_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a2bb2oi_1
X_06742_ _02647_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__buf_4
XFILLER_209_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._496_ AuI.pe._028_ AuI.pe._050_ AuI.pe._042_ AuI.pe._055_ AuI.pe._057_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._058_ sky130_fd_sc_hd__a221o_1
XMuI._4567_ MuI._0254_ MuI._0260_ MuI._0258_ vssd1 vssd1 vccd1 vccd1 MuI._0267_ sky130_fd_sc_hd__a21o_1
X_09461_ _02082_ _02084_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__or2b_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6306_ MuI._2077_ MuI._2120_ MuI._2179_ vssd1 vssd1 vccd1 vccd1 MuI._2180_ sky130_fd_sc_hd__a21bo_1
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3518_ MuI._0636_ MuI._0592_ MuI._0801_ MuI._0383_ vssd1 vssd1 vccd1 vccd1 MuI._1054_
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _06631_ _06630_ _04585_ _00048_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__and4_1
XFILLER_197_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4498_ MuI._0188_ MuI._0190_ vssd1 vssd1 vccd1 vccd1 MuI._0191_ sky130_fd_sc_hd__or2b_1
X_09392_ _01989_ _01985_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__or2b_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6237_ MuI._2860_ MuI._0515_ MuI._2008_ vssd1 vssd1 vccd1 vccd1 MuI._2104_ sky130_fd_sc_hd__and3_1
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12958__A1 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__B _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3449_ MuI.a_operand\[24\] MuI.b_operand\[24\] vssd1 vssd1 vccd1 vccd1 MuI._0295_
+ sky130_fd_sc_hd__nand2_1
X_08343_ _00958_ _00959_ _00960_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__o21bai_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6168_ MuI._0790_ MuI._2796_ vssd1 vssd1 vccd1 vccd1 MuI._2028_ sky130_fd_sc_hd__nand2_1
XFILLER_177_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3884__B MuI._2840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _00882_ _00889_ _00890_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__a21oi_1
XFILLER_193_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5119_ MuI.a_operand\[13\] MuI.a_operand\[12\] MuI._0017_ MuI._0018_ vssd1 vssd1
+ vccd1 vccd1 MuI._0874_ sky130_fd_sc_hd__and4_1
X_07225_ _02528_ _06525_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__nand2_1
XFILLER_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07021__A _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6099_ MuI._1950_ MuI._1951_ vssd1 vssd1 vccd1 vccd1 MuI._1952_ sky130_fd_sc_hd__nor2_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07156_ _06455_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__and2_1
XFILLER_180_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06860__A _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09874__C _06437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0989__A1 net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07087_ _04800_ _06284_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__and2_1
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13135__A1 _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout111 net59 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_6
Xfanout122 net39 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_6
Xfanout133 net12 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_4
XFILLER_102_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08787__A _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07691__A _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07989_ _00312_ _00603_ _00606_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__a21o_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09728_ _02348_ _02349_ _02365_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08314__A1 _00915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12459__D _05498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _02296_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__o21bai_1
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _05528_ _05538_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _00262_ _05262_ _04411_ _04210_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a31o_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4460__A1 MuI.a_operand\[20\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09130__B _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11621__A1 _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _04325_ _04337_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6170__B MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _03029_ _03027_ _03028_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__a21bo_1
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0930_ net20 AuI._0119_ AuI._0120_ vssd1 vssd1 vccd1 vccd1 AuI._0142_ sky130_fd_sc_hd__or3_1
XFILLER_184_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10707__D _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11483_ _04261_ _04263_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__xnor2_2
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__D _05101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12177__A2 _02736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13222_ _06128_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__nor2_1
X_10434_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0861_ AuI._0053_ net34 AuI._0080_ net106 vssd1 vssd1 vccd1 vccd1 AuI._0081_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_183_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06770__A _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11388__A _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _03055_ _03057_ _03058_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a21o_1
X_13153_ _06055_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__or2_1
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10723__C _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _04927_ _04928_ _04930_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a21o_1
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13084_ _03831_ _05467_ _05897_ _05894_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a31o_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _00345_ _04380_ _02982_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a22o_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10202__A_N _02259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ _04813_ _04814_ _04856_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__nor4_2
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._581__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1413_ AuI._0596_ AuI._0600_ vssd1 vssd1 vccd1 vccd1 AuI._0601_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5470_ MuI._1243_ MuI._1244_ MuI._1259_ vssd1 vssd1 vccd1 vccd1 MuI._1260_ sky130_fd_sc_hd__nand3_2
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1344_ AuI._0486_ AuI._0490_ AuI._0501_ AuI._0516_ vssd1 vssd1 vccd1 vccd1 AuI._0539_
+ sky130_fd_sc_hd__and4_1
XANTENNA__12012__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4421_ MuI.b_operand\[21\] MuI._3247_ MuI._3372_ MuI._2826_ vssd1 vssd1 vccd1
+ vccd1 MuI._0106_ sky130_fd_sc_hd__a22oi_1
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07106__A _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _05780_ _05781_ _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o21ai_1
XAuI._1275_ AuI._0420_ AuI._0465_ AuI._0474_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0475_
+ sky130_fd_sc_hd__a31o_1
XFILLER_207_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3688__C MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4352_ MuI._0029_ MuI._0030_ vssd1 vssd1 vccd1 vccd1 MuI._0031_ sky130_fd_sc_hd__nor2_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06945__A _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ _05359_ _05749_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a21bo_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4283_ MuI._3242_ MuI._3248_ MuI._3243_ vssd1 vssd1 vccd1 vccd1 MuI._3383_ sky130_fd_sc_hd__o21ba_1
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ _04607_ _02941_ _02731_ AuI.result\[10\] vssd1 vssd1 vccd1 vccd1 _04626_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6022_ MuI._1865_ MuI._1866_ vssd1 vssd1 vccd1 vccd1 MuI._1867_ sky130_fd_sc_hd__nor2_1
X_12799_ MuI.result\[19\] _02736_ _02944_ _05134_ _05678_ vssd1 vssd1 vccd1 vccd1
+ _05679_ sky130_fd_sc_hd__a221o_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07479__C _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6080__B MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__B _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07010_ _05531_ _05069_ _05144_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_1
XFILLER_162_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11729__C _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6855_ MuI._2672_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[22\] sky130_fd_sc_hd__nor2_1
XFILLER_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5424__B MuI._2875_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _03174_ _03971_ _01205_ _01207_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a22oi_1
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5806_ MuI._1595_ MuI._1596_ MuI._1627_ MuI._1628_ vssd1 vssd1 vccd1 vccd1 MuI._1630_
+ sky130_fd_sc_hd__o22a_1
XMuI._6786_ MuI._2505_ MuI._2563_ MuI._2559_ MuI._2567_ vssd1 vssd1 vccd1 vccd1 MuI._2708_
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07912_ _05370_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__buf_4
XMuI._3998_ MuI._3092_ MuI._3096_ MuI._3097_ vssd1 vssd1 vccd1 vccd1 MuI._3098_ sky130_fd_sc_hd__nand3_1
XANTENNA_AuI.pe._572__A2 AuI.pe._050_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08892_ _01357_ _01353_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__and2b_1
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5737_ MuI._1552_ MuI._1553_ vssd1 vssd1 vccd1 vccd1 MuI._1554_ sky130_fd_sc_hd__nor2_1
XANTENNA_AuI.pe._408__A AuI.pe.significand\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1396__A1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__A2 _05456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07843_ _03152_ _04638_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__nand2_1
XFILLER_112_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._617_ AuI.pe._162_ AuI.pe._163_ AuI.pe._166_ AuI.pe._169_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[13\] sky130_fd_sc_hd__o31a_1
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5668_ MuI._1476_ MuI._1477_ vssd1 vssd1 vccd1 vccd1 MuI._1478_ sky130_fd_sc_hd__nor2_1
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08757__D _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _00389_ _00390_ _00391_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__nand3_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6255__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4619_ MuI._0314_ MuI._0323_ vssd1 vssd1 vccd1 vccd1 MuI._0324_ sky130_fd_sc_hd__xor2_1
XAuI.pe._548_ AuI.pe.significand\[9\] vssd1 vssd1 vccd1 vccd1 AuI.pe._105_ sky130_fd_sc_hd__buf_2
XANTENNA__07016__A _05595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09513_ _02074_ _02086_ _02081_ _02085_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__o211a_1
XANTENNA__07676__A1_N _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5599_ MuI._1334_ MuI._1401_ vssd1 vssd1 vccd1 vccd1 MuI._1402_ sky130_fd_sc_hd__or2_1
X_06725_ net66 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__buf_4
XANTENNA_MuI._4056__A MuI._3154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._479_ AuI.pe._037_ AuI.pe._038_ AuI.pe._039_ AuI.pe._042_ AuI.pe._030_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._043_ sky130_fd_sc_hd__a32o_1
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ _02063_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nor2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06855__A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09375_ _01939_ _01942_ _01941_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12068__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10377__A _02431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08326_ _00908_ _00941_ _00942_ _00943_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__nand4_1
XFILLER_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08257_ net121 _04585_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__and2_1
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13356__A1 _04161_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07208_ _06498_ _06507_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a21bo_1
XFILLER_165_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08188_ _00804_ _00805_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__xnor2_2
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12742__D _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ _06439_ _06437_ _06432_ _06435_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11639__C _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13108__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10150_ _02827_ _05724_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nor2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _02216_ _03982_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__xnor2_4
XFILLER_181_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4892__C MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09125__B _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3484__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _03540_ _03542_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nand2_1
XANTENNA__12767__A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__A _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ _05594_ _02903_ _02925_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__mux2_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1060_ AuI._0269_ AuI._0270_ AuI._0189_ vssd1 vssd1 vccd1 vccd1 AuI._0271_ sky130_fd_sc_hd__mux2_1
XANTENNA__11842__A1 AuI.result\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A2 _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11842__B2 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06765__A _02894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12917__D _05649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ _05519_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10287__A _03798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _04190_ _04192_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__nand2_1
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12584_ _00290_ _00289_ _05509_ _03424_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nand4_2
XANTENNA__07299__C _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6186__A1 MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6186__B2 MuI._2814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ _04317_ _04318_ _04313_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._159_ FuI.a_operand\[29\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_144_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0913_ AuI._0130_ AuI._0131_ vssd1 vssd1 vccd1 vccd1 AuI._0132_ sky130_fd_sc_hd__or2_1
XFILLER_171_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _04241_ _04242_ _04243_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a21oi_1
XMuI._4970_ MuI._2693_ MuI._2638_ MuI._3362_ MuI._0100_ vssd1 vssd1 vccd1 vccd1 MuI._0710_
+ sky130_fd_sc_hd__and4_1
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07460__A2_N _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ _06110_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__xnor2_1
XAuI._0844_ net125 net109 vssd1 vssd1 vccd1 vccd1 AuI._0064_ sky130_fd_sc_hd__and2b_1
X_10417_ _00669_ _03114_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08223__B1 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11397_ FuI.Integer\[7\] _06056_ _04166_ _04167_ _04170_ vssd1 vssd1 vccd1 vccd1
+ _04171_ sky130_fd_sc_hd__a2111o_1
XFILLER_180_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3921_ MuI._0603_ MuI._2787_ MuI._2363_ MuI._2826_ vssd1 vssd1 vccd1 vccd1 MuI._3021_
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08219__A2_N _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _06036_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and2_1
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _03040_ _03041_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__nand2_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6640_ MuI._1238_ MuI._1458_ vssd1 vssd1 vccd1 vccd1 MuI._2547_ sky130_fd_sc_hd__and2b_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3852_ MuI._2937_ MuI._2951_ vssd1 vssd1 vccd1 vccd1 MuI._2952_ sky130_fd_sc_hd__xnor2_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _03744_ _05585_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a21o_1
X_10279_ _02964_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__xnor2_1
XMuI._6571_ MuI._2422_ MuI._2468_ MuI._2470_ MuI._2421_ vssd1 vssd1 vccd1 vccd1 MuI._2471_
+ sky130_fd_sc_hd__o211a_1
XMuI._3783_ MuI._0328_ MuI._2882_ vssd1 vssd1 vccd1 vccd1 MuI._2883_ sky130_fd_sc_hd__nand2_1
X_12018_ _04834_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand3_2
XMuI._5522_ MuI._1314_ MuI._1316_ vssd1 vssd1 vccd1 vccd1 MuI._1317_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09035__B _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._402_ AuI.pe.significand\[17\] AuI.pe.significand\[18\] AuI.pe.significand\[19\]
+ AuI.pe.significand\[20\] vssd1 vssd1 vccd1 vccd1 AuI.pe._369_ sky130_fd_sc_hd__or4_2
XMuI._5453_ MuI._1235_ MuI._1240_ vssd1 vssd1 vccd1 vccd1 MuI._1242_ sky130_fd_sc_hd__nand2_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1327_ AuI._0498_ AuI._0438_ AuI._0210_ vssd1 vssd1 vccd1 vccd1 AuI._0523_ sky130_fd_sc_hd__or3b_1
XFILLER_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4404_ MuI.a_operand\[7\] vssd1 vssd1 vccd1 vccd1 MuI._0088_ sky130_fd_sc_hd__clkbuf_4
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11581__A _02658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5384_ MuI._1156_ MuI._1163_ MuI._1165_ vssd1 vssd1 vccd1 vccd1 MuI._1166_ sky130_fd_sc_hd__and3_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07490_ _00056_ _00067_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__nand2_1
XFILLER_80_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1258_ AuI._0457_ AuI._0459_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[10\]
+ sky130_fd_sc_hd__xor2_2
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4335_ MuI._3305_ MuI._0012_ vssd1 vssd1 vccd1 vccd1 MuI._0013_ sky130_fd_sc_hd__xor2_2
XFILLER_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6091__A MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10197__A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1189_ net33 net65 AuI._0124_ vssd1 vssd1 vccd1 vccd1 AuI._0395_ sky130_fd_sc_hd__mux2_1
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4266_ MuI._3361_ MuI._3364_ MuI._3365_ vssd1 vssd1 vccd1 vccd1 MuI._3366_ sky130_fd_sc_hd__o21ba_1
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _02474_ _00082_ _00084_ _06564_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10628__C _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6005_ MuI._1847_ MuI._1848_ vssd1 vssd1 vccd1 vccd1 MuI._1849_ sky130_fd_sc_hd__xor2_2
XANTENNA__09201__D net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._490__A1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ _00727_ _00036_ _00059_ _00728_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__a22oi_1
XMuI._4197_ MuI._3285_ MuI._3294_ MuI._3295_ vssd1 vssd1 vccd1 vccd1 MuI._3297_ sky130_fd_sc_hd__or3_1
X_09091_ _01605_ _01606_ _01607_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a21oi_2
XFILLER_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08462__B1 _00090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10925__A _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08042_ _00658_ _00657_ _00656_ _00653_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__o211ai_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10644__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5292__A1_N MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08114__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _02651_ _02652_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__and2_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__B1_N _00664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6838_ MuI._2751_ vssd1 vssd1 vccd1 vccd1 MuI.result\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ _01549_ _01550_ _01560_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07953__B _02948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._545__A2 AuI.pe._070_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6769_ MuI._2588_ MuI._2597_ MuI._2601_ MuI._2688_ vssd1 vssd1 vccd1 vccd1 MuI._2689_
+ sky130_fd_sc_hd__and4_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08875_ _01448_ _01453_ _01447_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ net45 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__buf_6
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4663__A1 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07757_ _06460_ net128 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__and2_1
XANTENNA_MuI._5320__D MuI._0020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0914__A AuI._0132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11824__A1 _02669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06708_ net110 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__buf_4
XANTENNA__10627__A2 _04369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07688_ _00283_ _03971_ _00280_ _00282_ vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ _06519_ _06515_ net124 net123 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__and4_1
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5612__B1 MuI._0246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09896__A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ _01973_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__o21bai_1
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4959__A2_N MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08309_ _00918_ _00925_ _00926_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _01905_ _01902_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10260__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ _03938_ _03941_ _04086_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a211oi_4
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08305__A _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ _02442_ _04327_ _02744_ _06045_ FuI.Integer\[6\] vssd1 vssd1 vccd1 vccd1
+ _04014_ sky130_fd_sc_hd__a32o_1
XFILLER_107_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10202_ _02259_ _04057_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__and2b_1
X_11182_ _03936_ _03937_ _03921_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a21o_1
XFILLER_180_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _02795_ _02800_ _02805_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__and4b_1
XANTENNA_MuI._5999__B MuI._3156_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10064_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_input34_A a_operand[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07192__B1 _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07731__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0824__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1112_ AuI._0304_ AuI._0320_ AuI._0321_ AuI._0255_ vssd1 vssd1 vccd1 vccd1 AuI._0322_
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10618__A2 _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10966_ net60 _04380_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nand2_1
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10729__B _02229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1043_ net29 AuI._0138_ vssd1 vssd1 vccd1 vccd1 AuI._0255_ sky130_fd_sc_hd__xor2_1
X_12705_ _02970_ _04994_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nand2_1
XANTENNA__07495__A1 _06629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4424__A MuI.a_operand\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11291__A2 _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4120_ MuI._1274_ MuI._2787_ vssd1 vssd1 vccd1 vccd1 MuI._3220_ sky130_fd_sc_hd__nand2_1
X_10897_ _02388_ _05970_ _03630_ _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand4_2
XFILLER_204_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6342__C MuI._1494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _00299_ _00231_ _00385_ _00783_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__and4_1
XMuI._4051_ MuI._3089_ MuI._3150_ MuI._3070_ vssd1 vssd1 vccd1 vccd1 MuI._3151_ sky130_fd_sc_hd__or3_1
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._511__A AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12240__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._1296__B1 AuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12240__B2 _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _05427_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__xnor2_1
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11518_ _04298_ _04299_ _04136_ _04138_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__o211ai_2
XFILLER_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12498_ _04877_ _05352_ _05354_ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__a211o_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ _06620_ _03257_ _04224_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__nand4_1
XMuI._4953_ MuI._0602_ MuI._0690_ vssd1 vssd1 vccd1 vccd1 MuI._0692_ sky130_fd_sc_hd__or2_1
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0827_ net123 net107 vssd1 vssd1 vccd1 vccd1 AuI._0047_ sky130_fd_sc_hd__and2b_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3904_ MuI._2997_ MuI._3002_ MuI._3003_ vssd1 vssd1 vccd1 vccd1 MuI._3004_ sky130_fd_sc_hd__nand3_1
XFILLER_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08869__B _04907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4884_ MuI._2799_ MuI._2638_ MuI._0088_ MuI._2319_ vssd1 vssd1 vccd1 vccd1 MuI._0616_
+ sky130_fd_sc_hd__and4_1
XFILLER_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__xnor2_1
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _05316_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__clkbuf_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6623_ MuI._2526_ MuI._1433_ MuI._1434_ MuI._1444_ vssd1 vssd1 vccd1 vccd1 MuI._2529_
+ sky130_fd_sc_hd__nand4_1
XMuI._3835_ MuI._2927_ MuI._2934_ vssd1 vssd1 vccd1 vccd1 MuI._2935_ sky130_fd_sc_hd__xnor2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__A1 _00698_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6554_ MuI._2232_ MuI._2448_ vssd1 vssd1 vccd1 vccd1 MuI._2453_ sky130_fd_sc_hd__nor2_1
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3503__A MuI._0878_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3766_ MuI.b_operand\[7\] vssd1 vssd1 vccd1 vccd1 MuI._2866_ sky130_fd_sc_hd__buf_2
XFILLER_39_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08660_ _00983_ _00977_ _00982_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__nand3_1
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5505_ MuI._2892_ MuI._3185_ MuI._3371_ MuI._0110_ vssd1 vssd1 vccd1 vccd1 MuI._1299_
+ sky130_fd_sc_hd__and4_1
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6485_ MuI._2349_ MuI._2360_ vssd1 vssd1 vccd1 vccd1 MuI._2377_ sky130_fd_sc_hd__xnor2_1
X_07611_ _00225_ _00226_ _00227_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__a21o_1
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3697_ MuI._2539_ vssd1 vssd1 vccd1 vccd1 MuI._2797_ sky130_fd_sc_hd__buf_2
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08591_ _03174_ _04057_ _01158_ _01159_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_MuI._6814__A MuI.Exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5436_ MuI._1218_ MuI._1220_ MuI._1222_ vssd1 vssd1 vccd1 vccd1 MuI._1223_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07542_ _06475_ _05574_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__nand2_1
XANTENNA__12200__A _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10639__B _04197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5367_ MuI._2869_ MuI._0305_ MuI._0445_ MuI._2867_ vssd1 vssd1 vccd1 vccd1 MuI._1147_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__13092__B_N _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07473_ _00080_ _00087_ _00088_ _00090_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__and4bb_1
XMuI._4318_ MuI._3392_ MuI._3416_ MuI._3417_ vssd1 vssd1 vccd1 vccd1 MuI._3418_ sky130_fd_sc_hd__a21oi_2
XANTENNA_MuI._6252__C MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ _01696_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__and3_1
XFILLER_210_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5298_ MuI._0168_ MuI._3371_ MuI._0808_ MuI._0809_ vssd1 vssd1 vccd1 vccd1 MuI._1071_
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5070__A1 MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5070__B2 MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4249_ MuI.a_operand\[8\] vssd1 vssd1 vccd1 vccd1 MuI._3349_ sky130_fd_sc_hd__clkbuf_4
X_09143_ _01436_ _01618_ _01619_ _01620_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__and4b_1
XANTENNA__07948__B _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13031__A _04677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _01686_ _01687_ _01691_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__a21o_1
XFILLER_136_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__A1 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__C1 _05377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__B2 _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08025_ _00545_ _00560_ _00553_ _00559_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__a211o_1
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12534__A2 _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__B net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10390__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _01962_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__nor2_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08927_ _01537_ _01538_ _01544_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a21oi_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__D _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _06515_ _00032_ _04767_ net107 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__a22o_1
XANTENNA__10848__A2 _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4228__B MuI._2660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _00422_ _00426_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13247__B1 _06155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5050__D MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _01405_ _01406_ _03174_ _03884_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__and4bb_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _03536_ _03546_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__and3_1
XANTENNA__13206__A _02815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10549__B _03257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07204__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _03377_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5059__B MuI._3190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ _02820_ _06365_ _02814_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10682_ _03099_ _04961_ _06584_ _03056_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a22o_1
XFILLER_179_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _05270_ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__nor2_1
XFILLER_127_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08977__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5199__A1_N MuI._2895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08977__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ _05099_ _05104_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a211oi_4
XFILLER_154_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _00727_ _00421_ _00423_ _00728_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a22oi_1
X_12283_ _05120_ _05121_ _05035_ _04981_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__o211ai_2
XFILLER_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1661_ AuI._0014_ vssd1 vssd1 vccd1 vccd1 AuI.result\[27\] sky130_fd_sc_hd__clkbuf_1
X_11234_ _03994_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__and2b_1
XANTENNA_AuI._0819__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1592_ AuI._0259_ AuI._0764_ AuI._0765_ AuI._0760_ vssd1 vssd1 vccd1 vccd1 AuI.result\[12\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__and2_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10116_ _02786_ _02790_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__nand2_1
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11096_ _03840_ _03841_ _03843_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or4_1
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3620_ MuI._2143_ MuI._2165_ vssd1 vssd1 vccd1 vccd1 MuI._2176_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__B _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3551_ MuI._1362_ MuI._1406_ vssd1 vssd1 vccd1 vccd1 MuI._1417_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6270_ MuI._2126_ MuI._2139_ vssd1 vssd1 vccd1 vccd1 MuI._2140_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3482_ MuI._0636_ MuI._0537_ MuI._0394_ vssd1 vssd1 vccd1 vccd1 MuI._0658_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13116__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09313__B _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5221_ MuI._1813_ MuI._0420_ MuI._0985_ vssd1 vssd1 vccd1 vccd1 MuI._0986_ sky130_fd_sc_hd__and3_1
X_11998_ _03593_ _04961_ _06584_ _03539_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__a22o_1
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ _02764_ _03503_ _03683_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__o21a_1
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5152_ MuI._3223_ MuI.b_operand\[5\] vssd1 vssd1 vccd1 vccd1 MuI._0910_ sky130_fd_sc_hd__nand2_1
XFILLER_177_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1026_ net66 net34 AuI._0122_ vssd1 vssd1 vccd1 vccd1 AuI._0238_ sky130_fd_sc_hd__mux2_1
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4103_ MuI._2856_ MuI._2855_ vssd1 vssd1 vccd1 vccd1 MuI._3203_ sky130_fd_sc_hd__and2b_1
XANTENNA__06953__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3993__A MuI._2473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5083_ MuI._0821_ MuI._0820_ vssd1 vssd1 vccd1 vccd1 MuI._0835_ sky130_fd_sc_hd__and2b_1
XFILLER_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08871__C _06580_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _03315_ _05387_ _05397_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__a211o_1
XANTENNA__10475__A _03157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4034_ MuI._3131_ MuI._3132_ MuI._3127_ vssd1 vssd1 vccd1 vccd1 MuI._3134_ sky130_fd_sc_hd__a21o_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__A1 _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07640__B2 _03056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5985_ MuI._1806_ MuI._1807_ vssd1 vssd1 vccd1 vccd1 MuI._1827_ sky130_fd_sc_hd__nand2_1
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5713__A MuI._2852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4936_ MuI._0667_ MuI._0668_ vssd1 vssd1 vccd1 vccd1 MuI._0673_ sky130_fd_sc_hd__xnor2_1
X_09830_ _02393_ _02403_ _02406_ _02441_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._796_ AuI.pe._384_ AuI.pe._387_ vssd1 vssd1 vccd1 vccd1 AuI.pe._336_ sky130_fd_sc_hd__nand2_1
XMuI._4867_ MuI._0480_ MuI._0596_ vssd1 vssd1 vccd1 vccd1 MuI._0597_ sky130_fd_sc_hd__nor2_1
X_09761_ _06479_ net127 net126 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__and3_1
XFILLER_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06973_ _02140_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__clkbuf_2
XMuI._6606_ MuI._1766_ MuI._1815_ vssd1 vssd1 vccd1 vccd1 MuI._2510_ sky130_fd_sc_hd__and2b_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3818_ MuI.b_operand\[12\] vssd1 vssd1 vccd1 vccd1 MuI._2918_ sky130_fd_sc_hd__buf_2
X_08712_ _01328_ _01329_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__xor2_2
XMuI._4798_ MuI._0395_ MuI._0392_ MuI._0393_ vssd1 vssd1 vccd1 vccd1 MuI._0521_ sky130_fd_sc_hd__and3_1
XFILLER_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09692_ _02332_ _02331_ _02159_ _02147_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a211o_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3749_ MuI._2627_ vssd1 vssd1 vccd1 vccd1 MuI._2849_ sky130_fd_sc_hd__clkbuf_4
XMuI._6537_ MuI._2432_ MuI._2433_ vssd1 vssd1 vccd1 vccd1 MuI._2434_ sky130_fd_sc_hd__nor2_1
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08643_ _01259_ _01260_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__or2_1
XFILLER_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6468_ MuI._2354_ MuI._2356_ vssd1 vssd1 vccd1 vccd1 MuI._2358_ sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _01188_ _01190_ _01191_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__nor3_1
XANTENNA_MuI._4094__A2 MuI._2898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5419_ MuI._1148_ MuI._1147_ vssd1 vssd1 vccd1 vccd1 MuI._1204_ sky130_fd_sc_hd__nor2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6399_ MuI._2278_ MuI._2279_ MuI._2281_ vssd1 vssd1 vccd1 vccd1 MuI._2282_ sky130_fd_sc_hd__and3_1
X_07525_ _00121_ _00122_ _00141_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__nor3_4
XANTENNA__11255__A2 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08120__A2 _00735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ net123 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12584__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07387_ _00001_ _00003_ _06681_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a21o_1
XANTENNA__10385__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ _02905_ _02970_ _03884_ _03971_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__and4_1
XANTENNA__12755__A2 _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4511__B MuI._0182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09057_ _01626_ _01674_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12507__A2 _02738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _06491_ _05434_ _06466_ _06534_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__a22oi_2
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10832__B _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13180__A2 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1432__B1 AuI._0550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07395__B1 _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11191__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__B _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4884__D MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _02614_ _02609_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__nor2_1
XFILLER_131_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _02908_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nand2_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _04723_ _04733_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__and3_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11494__A2 _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12691__A1 _05559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _04505_ _04507_ _04368_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__a21oi_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _03517_ _03519_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__a21oi_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _04454_ _04459_ _04584_ _04586_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a211o_1
XFILLER_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08111__A2 _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ _03453_ _03455_ _03448_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a21o_1
XFILLER_186_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0821__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5585__A2 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4124__D MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _02921_ _06338_ _02824_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10665_ _00062_ _06525_ _06568_ _00063_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a22o_1
XANTENNA__10295__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _02795_ _05028_ _06629_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a21boi_1
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13384_ _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__or2_1
XFILLER_194_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10596_ _02259_ _04068_ _02743_ _06045_ FuI.Integer\[2\] vssd1 vssd1 vccd1 vccd1
+ _03309_ sky130_fd_sc_hd__a32o_1
XFILLER_126_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12335_ _05178_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nand2_1
XFILLER_182_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12266_ _05103_ _05104_ _05093_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5770_ MuI._1581_ MuI._1583_ MuI._1588_ vssd1 vssd1 vccd1 vccd1 MuI._1590_ sky130_fd_sc_hd__o21bai_1
X_11217_ _03970_ _03972_ _03975_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a21o_1
XAuI._1644_ AuI.exp_a AuI._0710_ AuI.operand_a\[24\] vssd1 vssd1 vccd1 vccd1 AuI._0001_
+ sky130_fd_sc_hd__a21oi_1
X_12197_ _02935_ _05029_ _05030_ _02732_ AuI.result\[14\] vssd1 vssd1 vccd1 vccd1
+ _05031_ sky130_fd_sc_hd__a32o_1
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 ALU_Output[10] sky130_fd_sc_hd__buf_2
XANTENNA__12015__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6298__B1 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._650_ AuI.pe._378_ AuI.pe._002_ AuI.pe._053_ AuI.pe.significand\[12\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._200_ sky130_fd_sc_hd__a22o_1
XMuI._4721_ MuI._0433_ MuI._0435_ vssd1 vssd1 vccd1 vccd1 MuI._0436_ sky130_fd_sc_hd__nand2_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 ALU_Output[20] sky130_fd_sc_hd__buf_2
XFILLER_123_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 ALU_Output[30] sky130_fd_sc_hd__buf_2
XFILLER_150_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11148_ _03774_ _03776_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__o211ai_4
XAuI._1575_ AuI._0693_ AuI._0746_ AuI._0750_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0751_
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4652_ MuI._0349_ MuI._0357_ MuI._0359_ vssd1 vssd1 vccd1 vccd1 MuI._0360_ sky130_fd_sc_hd__a21oi_1
XAuI.pe._581_ AuI.pe._102_ AuI.pe._050_ AuI.pe._079_ AuI.pe._063_ AuI.pe._135_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._136_ sky130_fd_sc_hd__a221o_1
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11079_ _03824_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__xnor2_4
XMuI._3603_ MuI._1923_ MuI._1956_ MuI._1978_ vssd1 vssd1 vccd1 vccd1 MuI._1989_ sky130_fd_sc_hd__o21a_1
XANTENNA__06948__A _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3520__A1 MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__B1 _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4583_ MuI._0279_ MuI._0277_ vssd1 vssd1 vccd1 vccd1 MuI._0285_ sky130_fd_sc_hd__xor2_1
XFILLER_209_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6322_ MuI._2146_ MuI._2148_ MuI._2196_ vssd1 vssd1 vccd1 vccd1 MuI._2197_ sky130_fd_sc_hd__o21ai_1
XMuI._3534_ MuI._1131_ MuI._1219_ vssd1 vssd1 vccd1 vccd1 MuI._1230_ sky130_fd_sc_hd__nand2_1
XFILLER_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4713__A2_N MuI._3247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__D _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__C _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10189__B _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6253_ MuI._0614_ MuI._3091_ MuI._2849_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._2122_
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3465_ MuI._0460_ vssd1 vssd1 vccd1 vccd1 MuI._0471_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09978__B _02637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5204_ MuI._0864_ MuI._0858_ MuI._0863_ vssd1 vssd1 vccd1 vccd1 MuI._0968_ sky130_fd_sc_hd__a21o_1
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6184_ MuI._2817_ MuI._3091_ vssd1 vssd1 vccd1 vccd1 MuI._2046_ sky130_fd_sc_hd__nand2_1
X_07310_ net9 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06683__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08290_ _00874_ _00905_ _00906_ _00907_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__a211o_1
XFILLER_189_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5135_ MuI._0887_ MuI._0891_ vssd1 vssd1 vccd1 vccd1 MuI._0892_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1009_ AuI._0190_ AuI._0191_ AuI._0220_ vssd1 vssd1 vccd1 vccd1 AuI._0221_ sky130_fd_sc_hd__or3b_1
X_07241_ _06539_ _06540_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__nand3_1
XANTENNA__12835__D _05574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4612__A MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5066_ MuI._2853_ MuI._2854_ MuI.a_operand\[4\] MuI.a_operand\[3\] vssd1 vssd1
+ vccd1 vccd1 MuI._0816_ sky130_fd_sc_hd__and4_1
X_07172_ _06465_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nand3_1
XFILLER_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4017_ MuI._3115_ MuI._3116_ vssd1 vssd1 vccd1 vccd1 MuI._3117_ sky130_fd_sc_hd__xnor2_2
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07945__C _00105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4985__C MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5968_ MuI._1806_ MuI._1807_ vssd1 vssd1 vccd1 vccd1 MuI._1808_ sky130_fd_sc_hd__xnor2_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6258__B MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4919_ MuI._0613_ MuI._0653_ vssd1 vssd1 vccd1 vccd1 MuI._0654_ sky130_fd_sc_hd__nand2_1
X_09813_ _02459_ _02460_ _02463_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__and3_1
XFILLER_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07019__A _05627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5899_ MuI._1729_ MuI._1730_ MuI._1679_ MuI._1720_ vssd1 vssd1 vccd1 vccd1 MuI._1732_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_87_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._779_ AuI.pe._399_ AuI.pe._078_ vssd1 vssd1 vccd1 vccd1 AuI.pe._320_ sky130_fd_sc_hd__or2_1
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09744_ _02287_ _02315_ _02314_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__and3_1
XFILLER_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06956_ net133 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__buf_4
XANTENNA__06858__A _03895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3898__A MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09675_ _02269_ _02316_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or2_1
XANTENNA__11476__A2 _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ _04208_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[4\] sky130_fd_sc_hd__clkbuf_2
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A2 _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08626_ _01091_ _01093_ _01104_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__nor3_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08557_ _00874_ _00902_ _00903_ _00904_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__and4_1
XANTENNA__08629__B1 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0922__A AuI._0136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12976__A2 _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07508_ _00124_ _00125_ _04445_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__and3_1
XFILLER_196_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08488_ _00882_ _00888_ _00887_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__a21o_1
XFILLER_211_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07439_ _06600_ _06609_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__nor2_1
XFILLER_211_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11004__A _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _06429_ _04197_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nand2_1
XFILLER_183_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5319__A2 MuI._3262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _01724_ _01725_ _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a21o_1
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07604__A1 _00221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _03074_ _03075_ _03070_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__a21o_1
XFILLER_124_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _04947_ _04948_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__xor2_2
XFILLER_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5353__A MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ _04612_ _04613_ _04759_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or3_1
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6168__B MuI._2796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _02894_ _00046_ _00412_ _00530_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__nand4_1
XFILLER_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1360_ AuI._0528_ AuI._0534_ AuI._0545_ AuI._0553_ vssd1 vssd1 vccd1 vccd1 AuI._0554_
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06768__A _02927_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _01962_ _02640_ _05757_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__and3_1
XANTENNA__12664__A1 _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1291_ AuI._0487_ AuI._0488_ AuI._0489_ vssd1 vssd1 vccd1 vccd1 AuI._0490_ sky130_fd_sc_hd__or3_2
XANTENNA_MuI._6184__A MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11904_ _04705_ _04706_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a21oi_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ FuI.Integer\[20\] _06056_ _04642_ _05209_ _05769_ vssd1 vssd1 vccd1 vccd1
+ _05770_ sky130_fd_sc_hd__a221o_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11835_ _02944_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__clkbuf_4
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09817__C1 _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07599__A _00028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12967__A2 _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _04565_ _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__xor2_4
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10717_ _03435_ _03436_ _03418_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a21o_1
X_11697_ _04493_ _02891_ _02928_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__mux2_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13436_ _05788_ _04642_ _06346_ _03680_ _06350_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a221o_1
X_10648_ _03361_ _03362_ _03358_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a21o_1
XFILLER_155_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _06231_ _06234_ _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__o21a_1
XFILLER_155_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ _03135_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__xnor2_2
XFILLER_127_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6871_ MuI._2735_ MuI._2771_ MuI._2761_ vssd1 vssd1 vccd1 vccd1 MuI.result\[27\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_115_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12318_ _03335_ _05520_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__nand2_1
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _02679_ _06207_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nand2_2
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5822_ MuI._1476_ MuI._1636_ MuI._1635_ vssd1 vssd1 vccd1 vccd1 MuI._1647_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09348__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12959__A1_N _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09348__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12249_ _04947_ _04948_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__and2_1
XAuI.pe._702_ AuI.pe._385_ AuI.pe._022_ AuI.pe._247_ AuI.pe._248_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._249_ sky130_fd_sc_hd__a211o_1
XFILLER_123_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5753_ MuI._1569_ MuI._1570_ vssd1 vssd1 vccd1 vccd1 MuI._1572_ sky130_fd_sc_hd__nand2_1
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1627_ AuI.pe.Significand\[19\] AuI._0695_ AuI._0760_ AuI._0793_ vssd1 vssd1
+ vccd1 vccd1 AuI.result\[19\] sky130_fd_sc_hd__o211a_1
XFILLER_111_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._633_ AuI.pe._170_ AuI.pe._167_ vssd1 vssd1 vccd1 vccd1 AuI.pe._184_ sky130_fd_sc_hd__or2_1
XMuI._4704_ MuI._0285_ MuI._0417_ vssd1 vssd1 vccd1 vccd1 MuI._0418_ sky130_fd_sc_hd__nand2_1
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ _03378_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__buf_4
XMuI._5684_ MuI._2583_ MuI._0112_ vssd1 vssd1 vccd1 vccd1 MuI._1496_ sky130_fd_sc_hd__nand2_1
XANTENNA__07781__B _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1558_ AuI._0645_ AuI._0651_ AuI._0663_ AuI._0666_ vssd1 vssd1 vccd1 vccd1 AuI._0737_
+ sky130_fd_sc_hd__and4_1
X_07790_ _00373_ _00185_ _00406_ _00407_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__o211ai_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._564_ AuI.pe.significand\[15\] vssd1 vssd1 vccd1 vccd1 AuI.pe._120_ sky130_fd_sc_hd__buf_2
XMuI._4635_ MuI.a_operand\[18\] MuI.a_operand\[17\] MuI._2884_ MuI._2880_ vssd1 vssd1
+ vccd1 vccd1 MuI._0342_ sky130_fd_sc_hd__and4_1
XFILLER_83_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4029__D MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ net38 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1489_ AuI._0674_ AuI._0670_ vssd1 vssd1 vccd1 vccd1 AuI._0675_ sky130_fd_sc_hd__nor2_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4566_ MuI._0264_ MuI._0265_ vssd1 vssd1 vccd1 vccd1 MuI._0266_ sky130_fd_sc_hd__xnor2_1
XAuI.pe._495_ AuI.pe._045_ AuI.pe._023_ AuI.pe._027_ AuI.pe._056_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._057_ sky130_fd_sc_hd__a22o_1
XANTENNA_AuI._0900__A_N net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _02083_ _02080_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6305_ MuI._0625_ MuI._2077_ MuI._3091_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._2179_
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3517_ MuI._1032_ vssd1 vssd1 vccd1 vccd1 MuI._1043_ sky130_fd_sc_hd__buf_2
XFILLER_52_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08411_ _02851_ _04531_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__nand2_1
XMuI._4497_ MuI._0052_ MuI._0189_ vssd1 vssd1 vccd1 vccd1 MuI._0190_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _01982_ _01984_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__or2b_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6236_ MuI._2073_ MuI._2074_ MuI._2101_ vssd1 vssd1 vccd1 vccd1 MuI._2103_ sky130_fd_sc_hd__a21o_1
XMuI._3448_ MuI.a_operand\[25\] MuI.b_operand\[25\] vssd1 vssd1 vccd1 vccd1 MuI._0284_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12958__A2 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _06469_ _02194_ net18 net19 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__and4_1
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6167_ MuI._2018_ MuI._2025_ MuI._2024_ vssd1 vssd1 vccd1 vccd1 MuI._2027_ sky130_fd_sc_hd__a21o_1
XANTENNA__07302__A _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ _00882_ _00889_ _00890_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._3884__C MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4342__A MuI._0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5118_ MuI._0477_ MuI._0378_ vssd1 vssd1 vccd1 vccd1 MuI._0873_ sky130_fd_sc_hd__nand2_1
XFILLER_165_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08117__B _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6098_ MuI._0372_ MuI._0625_ MuI._2797_ MuI._2789_ vssd1 vssd1 vccd1 vccd1 MuI._1951_
+ sky130_fd_sc_hd__and4_1
X_07224_ _05176_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__buf_4
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5049_ MuI._0085_ MuI._3306_ MuI._2881_ MuI._2341_ vssd1 vssd1 vccd1 vccd1 MuI._0797_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__09587__A1 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07155_ _03561_ _03615_ _03895_ _03993_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__and4_2
XFILLER_180_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09874__D _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07086_ _06336_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[12\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11478__B _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__C _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5173__A MuI._2853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13135__A2 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout112 net56 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_4
Xfanout123 net33 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_4
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__B _01206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07691__B _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5485__A1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07988_ _03324_ _04046_ _00604_ _00605_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__a31o_1
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09727_ _02370_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__xnor2_1
X_06939_ _04767_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_MuI._4517__A MuI._2799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09658_ _06469_ _00150_ net123 _00089_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__and4_1
XFILLER_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08609_ _01027_ _01028_ _01033_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__a21o_1
XFILLER_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09589_ _02179_ _02178_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__and2b_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11620_ _00132_ _05316_ _05380_ _00133_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__a22o_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__C _06666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13214__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08078__A1 _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4460__A2 MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08308__A _00596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07212__A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _02772_ _02889_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nand2_1
XANTENNA__07825__A1 _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07825__B2 _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11621__A2 _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6170__C MuI._2802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _03205_ _03203_ _03204_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nand3_1
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ _03722_ _04596_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__and2_1
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ _06125_ _06127_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nor2_1
X_10433_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__clkbuf_4
XAuI._0860_ net35 vssd1 vssd1 vccd1 vccd1 AuI._0080_ sky130_fd_sc_hd__inv_2
XFILLER_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A b_operand[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _06015_ _05971_ _06054_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__and3_1
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10364_ _03055_ _03057_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nand3_1
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _04927_ _04928_ _04930_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__and3_1
XFILLER_112_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10723__D _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _05908_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10295_ _02983_ _02984_ _00093_ _04520_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__nand4_2
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08978__A _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12034_ _04853_ _04855_ _04815_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12885__A1 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1412_ AuI._0597_ AuI._0598_ AuI.pe.significand\[24\] vssd1 vssd1 vccd1 vccd1
+ AuI._0600_ sky130_fd_sc_hd__o21a_1
XFILLER_78_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1343_ AuI._0518_ AuI._0524_ AuI._0537_ vssd1 vssd1 vccd1 vccd1 AuI._0538_ sky130_fd_sc_hd__o21ai_1
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4427__A MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4420_ MuI._0098_ MuI._0104_ vssd1 vssd1 vccd1 vccd1 MuI._0105_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12012__B _03271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09502__A1 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XAuI._1274_ AuI._0473_ vssd1 vssd1 vccd1 vccd1 AuI._0474_ sky130_fd_sc_hd__inv_2
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12936_ _05784_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__xor2_1
XFILLER_206_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4351_ MuI._0790_ MuI._1021_ MuI._2886_ MuI._2882_ vssd1 vssd1 vccd1 vccd1 MuI._0030_
+ sky130_fd_sc_hd__and4_1
XANTENNA_MuI._3688__D MuI._2773_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._514__A AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _05567_ _05568_ _05667_ _05750_ _05666_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a311oi_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4282_ MuI._3340_ MuI._3380_ MuI._3381_ vssd1 vssd1 vccd1 vccd1 MuI._3382_ sky130_fd_sc_hd__o21bai_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ _02860_ _04624_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6021_ MuI._1153_ MuI._2914_ MuI._2594_ MuI._0746_ vssd1 vssd1 vccd1 vccd1 MuI._1866_
+ sky130_fd_sc_hd__a22oi_1
X_12798_ _02720_ _02868_ _03973_ _02742_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ _04547_ _04548_ _04398_ _04419_ vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__o211a_1
XFILLER_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4162__A MuI.b_operand\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07479__D _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ _06330_ _06331_ _03133_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__o21a_1
XFILLER_190_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._0989_ net51 net19 AuI._0123_ vssd1 vssd1 vccd1 vccd1 AuI._0201_ sky130_fd_sc_hd__mux2_1
XANTENNA__11729__D _05316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6854_ MuI._2674_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[21\] sky130_fd_sc_hd__nor2_1
XFILLER_142_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._557__B1 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ _03239_ _03906_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__nand2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5805_ MuI._1595_ MuI._1596_ MuI._1627_ MuI._1628_ vssd1 vssd1 vccd1 vccd1 MuI._1629_
+ sky130_fd_sc_hd__nor4_2
X_07911_ _02377_ _06561_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__nand2_1
XFILLER_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6785_ MuI._2577_ MuI._2706_ vssd1 vssd1 vccd1 vccd1 MuI._2707_ sky130_fd_sc_hd__nor2_1
XMuI._3997_ MuI._3094_ MuI._3095_ MuI._3093_ vssd1 vssd1 vccd1 vccd1 MuI._3097_ sky130_fd_sc_hd__a21bo_1
X_08891_ _01507_ _01506_ _01481_ _01470_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o211a_1
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5736_ MuI._1550_ MuI._1551_ MuI._0990_ vssd1 vssd1 vccd1 vccd1 MuI._1553_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._408__B AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07842_ _00458_ _00459_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__xor2_2
XFILLER_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._616_ AuI.pe._167_ AuI.pe._168_ AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 AuI.pe._169_
+ sky130_fd_sc_hd__a21o_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5667_ MuI._1009_ MuI._1466_ MuI._1475_ vssd1 vssd1 vccd1 vccd1 MuI._1477_ sky130_fd_sc_hd__and3_1
X_07773_ _00380_ _00381_ _00388_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__a21o_1
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._547_ AuI.pe._094_ AuI.pe._100_ AuI.pe._104_ vssd1 vssd1 vccd1 vccd1 AuI.pe.Significand\[8\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4618_ MuI._0319_ MuI._0322_ vssd1 vssd1 vccd1 vccd1 MuI._0323_ sky130_fd_sc_hd__xnor2_1
X_09512_ _02136_ _02137_ _02120_ _02123_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__o211a_1
X_06724_ _02453_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_25_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5598_ MuI._1370_ MuI._1374_ MuI._1376_ MuI._1400_ vssd1 vssd1 vccd1 vccd1 MuI._1401_
+ sky130_fd_sc_hd__nand4_1
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._478_ AuI.pe._041_ vssd1 vssd1 vccd1 vccd1 AuI.pe._042_ sky130_fd_sc_hd__clkbuf_4
XMuI._4549_ MuI._0246_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._0247_ sky130_fd_sc_hd__nand2_1
X_09443_ _02063_ _02065_ net122 _06436_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and4bb_1
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _01981_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__nand3_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10377__B _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6219_ MuI._2041_ MuI._2075_ MuI._2082_ vssd1 vssd1 vccd1 vccd1 MuI._2084_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07032__A _05767_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _00907_ _00906_ _00905_ _00874_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__o211ai_2
XFILLER_178_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4072__A MuI._3160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12800__B2 _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10811__B1 _00040_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ _00849_ _00871_ _00872_ _00873_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__o211ai_4
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06871__A _04035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ _06486_ _06497_ _06487_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__nand3_1
XFILLER_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08187_ _00439_ _00477_ _00438_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a21boi_1
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07138_ net58 vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__buf_2
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13108__A2 _05999_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _06160_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11119__B2 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10080_ _02751_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__buf_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13209__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10195__B_N _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4892__D MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12619__A1 _03315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _03719_ _03720_ _03716_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a21o_1
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12767__B _05262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ _02856_ _05487_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a21o_1
XANTENNA__09422__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__A2 _02732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12652_ net60 _05262_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__and2_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__B _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ _04389_ _04390_ _04386_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__a21o_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5078__A MuI._2836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _00289_ _00398_ _03424_ _03378_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__a22o_1
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07299__D _04896_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11534_ _03657_ _04006_ _03832_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6186__A2 MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06781__A _03067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._158_ FuI.a_operand\[28\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[28\] sky130_fd_sc_hd__clkbuf_1
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0912_ AuI._0128_ AuI._0129_ AuI._0104_ vssd1 vssd1 vccd1 vccd1 AuI._0131_ sky130_fd_sc_hd__a21oi_1
XFILLER_172_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11465_ _04241_ _04242_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__and3_1
XFILLER_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._089_ FuI._051_ vssd1 vssd1 vccd1 vccd1 FuI._018_ sky130_fd_sc_hd__clkbuf_1
X_13204_ _03680_ _05777_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__nand2_1
XFILLER_99_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _00807_ _00808_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__nor2_1
XANTENNA__08223__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0843_ net110 AuI._0062_ net111 AuI._0057_ vssd1 vssd1 vccd1 vccd1 AuI._0063_
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ _04467_ _03675_ _02938_ AuI.result\[7\] _04169_ vssd1 vssd1 vccd1 vccd1 _04170_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__08223__B2 _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3920_ MuI._3018_ MuI._3019_ vssd1 vssd1 vccd1 vccd1 MuI._3020_ sky130_fd_sc_hd__nand2_1
XFILLER_180_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _03507_ _05981_ _05869_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__a31oi_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10347_ _03038_ _03039_ _03006_ _00768_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__o211ai_1
XFILLER_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3851_ MuI._2949_ MuI._2950_ vssd1 vssd1 vccd1 vccd1 MuI._2951_ sky130_fd_sc_hd__or2_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _03744_ _05585_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__nand3_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10278_ _02965_ _04186_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__nand2_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5541__A MuI._2966_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3782_ MuI._2881_ vssd1 vssd1 vccd1 vccd1 MuI._2882_ sky130_fd_sc_hd__buf_2
XMuI._6570_ MuI._2445_ MuI._2469_ vssd1 vssd1 vccd1 vccd1 MuI._2470_ sky130_fd_sc_hd__nand2_1
X_12017_ _00283_ _00423_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nand4_2
XFILLER_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5521_ MuI._1266_ MuI._1315_ vssd1 vssd1 vccd1 vccd1 MuI._1316_ sky130_fd_sc_hd__or2_1
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._401_ AuI.pe.significand\[21\] AuI.pe.significand\[23\] AuI.pe.significand\[22\]
+ AuI.pe.significand\[24\] vssd1 vssd1 vccd1 vccd1 AuI.pe._368_ sky130_fd_sc_hd__or4b_4
XFILLER_54_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5452_ MuI._1234_ MuI._1229_ MuI._1233_ vssd1 vssd1 vccd1 vccd1 MuI._1240_ sky130_fd_sc_hd__or3_1
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1326_ AuI._0513_ AuI._0522_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[15\]
+ sky130_fd_sc_hd__xnor2_4
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__B1 _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__A net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4403_ MuI._1296_ MuI.b_operand\[15\] MuI._2341_ MuI._0085_ vssd1 vssd1 vccd1
+ vccd1 MuI._0087_ sky130_fd_sc_hd__and4_1
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5383_ MuI._1154_ MuI._1155_ MuI._1139_ MuI._1152_ vssd1 vssd1 vccd1 vccd1 MuI._1165_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11581__B net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _03669_ _05520_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__nand2_1
XAuI._1257_ AuI._0434_ AuI._0447_ AuI._0458_ vssd1 vssd1 vccd1 vccd1 AuI._0459_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12192__A1_N _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4334_ MuI._3387_ MuI._0009_ MuI._0011_ vssd1 vssd1 vccd1 vccd1 MuI._0012_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13035__A1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13035__B2 _05338_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1188_ AuI._0367_ AuI._0382_ AuI._0392_ vssd1 vssd1 vccd1 vccd1 AuI._0394_ sky130_fd_sc_hd__nand3_1
XANTENNA_MuI._6091__B MuI._2813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4265_ MuI.b_operand\[19\] MuI._2811_ MuI._2374_ MuI._2319_ vssd1 vssd1 vccd1
+ vccd1 MuI._3365_ sky130_fd_sc_hd__and4_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10628__D _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6004_ MuI._3113_ MuI._3116_ MuI._3114_ vssd1 vssd1 vccd1 vccd1 MuI._1848_ sky130_fd_sc_hd__o21ba_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ _00299_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__buf_4
XMuI._4196_ MuI._3285_ MuI._3294_ MuI._3295_ vssd1 vssd1 vccd1 vccd1 MuI._3296_ sky130_fd_sc_hd__o21ai_1
X_09090_ _01696_ _01706_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__nand3_1
XANTENNA__08462__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06691__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ _00653_ _00656_ _00657_ _00658_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__a211o_1
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11349__A1 _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10644__C _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _02650_ _02655_ _02656_ _02657_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o211ai_2
XANTENNA_AuI._0813__A1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6837_ MuI._2690_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2751_ sky130_fd_sc_hd__and2b_1
XFILLER_115_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08943_ _01551_ _01552_ _01559_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__nand3_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07953__C _00098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__A _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6768_ MuI._2686_ MuI._2617_ vssd1 vssd1 vccd1 vccd1 MuI._2688_ sky130_fd_sc_hd__nor2_1
XFILLER_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11475__C _00033_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _01485_ _01486_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__nand3_1
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5719_ MuI._1524_ MuI._1532_ MuI._1533_ vssd1 vssd1 vccd1 vccd1 MuI._1534_ sky130_fd_sc_hd__nand3_1
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ _02840_ _00197_ _00199_ _00010_ _05123_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__a32o_1
XANTENNA__07027__A _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6699_ MuI._2505_ MuI._2599_ MuI._2610_ MuI._2611_ vssd1 vssd1 vccd1 vccd1 MuI._2612_
+ sky130_fd_sc_hd__a211o_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07756_ _06534_ _02205_ _00153_ net29 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__nand4_1
XANTENNA__06866__A _03982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4663__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06707_ _02270_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11824__A2 _02724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07687_ _00300_ _00304_ vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__nor2_1
XFILLER_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09426_ _06663_ _04176_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__nand2_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5612__A1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4514__B MuI._0208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09357_ _02096_ _02194_ net7 net8 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__and4_1
XANTENNA__09896__B _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0930__A net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08308_ _00596_ _00919_ _00924_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__and3_1
XFILLER_138_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09288_ _01902_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__and2b_1
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10260__B2 _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08239_ _00851_ _00856_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__and2_1
XFILLER_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08305__B _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ MuI.result\[6\] _02739_ _02719_ _04391_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_
+ sky130_fd_sc_hd__a221o_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__A2_N _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ _02302_ _04122_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__and2b_1
XFILLER_107_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ _03921_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand3_2
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _02806_ _02807_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__nor2b_2
XANTENNA__11760__B2 _04854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _02129_ _02064_ _02031_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__and3_2
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input27_A a_operand[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__A1 _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07192__B2 _06492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09469__B1 _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06776__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09152__A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1111_ AuI._0304_ AuI._0320_ vssd1 vssd1 vccd1 vccd1 AuI._0321_ sky130_fd_sc_hd__nand2_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10298__A _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__xor2_4
XFILLER_189_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12704_ _02623_ _05573_ _05576_ _03314_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__o211a_2
XANTENNA__10729__C _03247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1042_ AuI._0139_ AuI._0253_ vssd1 vssd1 vccd1 vccd1 AuI._0254_ sky130_fd_sc_hd__nor2_1
X_10896_ _03628_ _03629_ _03621_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__a21o_1
XFILLER_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6342__D MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12635_ _01146_ _03247_ _05820_ _03228_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a22oi_1
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4050_ MuI._3062_ MuI._3063_ vssd1 vssd1 vccd1 vccd1 MuI._3150_ sky130_fd_sc_hd__nor2_1
XANTENNA__13303__A2_N _02727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4143__C MuI._2330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _03658_ _05262_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__nand2_1
XFILLER_200_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12240__A2 _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5367__B1 MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11517_ _04136_ _04138_ _04298_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a211o_1
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4440__A MuI._0075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ _05242_ _05239_ _05238_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__o21ba_1
XFILLER_184_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output95_A net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _02593_ _02658_ _03082_ _00789_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nand4_2
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4952_ MuI._0599_ MuI._0601_ vssd1 vssd1 vccd1 vccd1 MuI._0690_ sky130_fd_sc_hd__nor2_1
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0826_ AuI._0037_ AuI._0043_ AuI._0045_ AuI._0041_ AuI._0040_ vssd1 vssd1 vccd1
+ vccd1 AuI._0046_ sky130_fd_sc_hd__a32o_1
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10761__A _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _03859_ _04000_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__o21ba_1
XFILLER_180_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3903_ MuI._2999_ MuI._3001_ MuI._2998_ vssd1 vssd1 vccd1 vccd1 MuI._3003_ sky130_fd_sc_hd__a21bo_1
XFILLER_180_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07955__B1 _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _03669_ _05713_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__nand2_1
XMuI._4883_ MuI._0528_ MuI._0612_ MuI._0611_ MuI._0588_ vssd1 vssd1 vccd1 vccd1 MuI._0615_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_113_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6622_ MuI._2526_ MuI._1445_ vssd1 vssd1 vccd1 vccd1 MuI._2527_ sky130_fd_sc_hd__or2b_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3834_ MuI._2928_ MuI._2933_ vssd1 vssd1 vccd1 vccd1 MuI._2934_ sky130_fd_sc_hd__xor2_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _03497_ _05842_ _05941_ _05943_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a22oi_1
XFILLER_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10306__A2 _00702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6553_ MuI._2205_ MuI._2206_ MuI._2450_ vssd1 vssd1 vccd1 vccd1 MuI._2452_ sky130_fd_sc_hd__o21ai_1
XMuI._3765_ MuI._2858_ MuI._2864_ vssd1 vssd1 vccd1 vccd1 MuI._2865_ sky130_fd_sc_hd__nand2_2
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5504_ MuI._2882_ MuI._0305_ MuI._0445_ MuI._2886_ vssd1 vssd1 vccd1 vccd1 MuI._1298_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07610_ _00225_ _00226_ _00227_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__nand3_1
XMuI._6484_ MuI._2372_ MuI._2375_ vssd1 vssd1 vccd1 vccd1 MuI._2376_ sky130_fd_sc_hd__or2b_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3696_ MuI.b_operand\[14\] vssd1 vssd1 vccd1 vccd1 MuI._2796_ sky130_fd_sc_hd__clkbuf_4
X_08590_ _03174_ _03971_ _01205_ _01207_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__and4_1
XFILLER_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5435_ MuI._1063_ MuI._1221_ vssd1 vssd1 vccd1 vccd1 MuI._1222_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._6814__B MuI._2731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1309_ AuI._0437_ AuI._0502_ AuI._0505_ AuI._0506_ vssd1 vssd1 vccd1 vccd1 AuI._0507_
+ sky130_fd_sc_hd__and4_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07541_ _00155_ _00157_ _00156_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a21o_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12200__B _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5366_ MuI._2871_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._1146_ sky130_fd_sc_hd__nand2_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ _00089_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__buf_4
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4317_ MuI._3413_ MuI._3415_ vssd1 vssd1 vccd1 vccd1 MuI._3417_ sky130_fd_sc_hd__and2_1
X_09211_ _01696_ _01707_ _01706_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5297_ MuI._2967_ MuI._2830_ MuI._1068_ MuI._1069_ vssd1 vssd1 vccd1 vccd1 MuI._1070_
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4248_ MuI._3345_ MuI._3347_ vssd1 vssd1 vccd1 vccd1 MuI._3348_ sky130_fd_sc_hd__or2b_1
X_09142_ _01618_ _01619_ _01759_ _01436_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13312__A _02830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4179_ MuI._3168_ MuI._3169_ vssd1 vssd1 vccd1 vccd1 MuI._3279_ sky130_fd_sc_hd__xnor2_2
XFILLER_163_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07310__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _01688_ _01689_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__o21bai_1
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10793__A2 _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08024_ _00640_ _00639_ _00638_ _00635_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__o211a_1
XANTENNA_MuI._4030__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13192__B1 _02713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11767__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__C _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _01844_ _02585_ _02037_ _01960_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__or4bb_1
XFILLER_131_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10390__B _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__A1_N _00444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _01539_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ net107 net66 net8 _04767_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__and4_1
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0925__A AuI._0116_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4228__C MuI._2844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07808_ _00424_ _00425_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__nor2_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _03110_ _06437_ _04046_ _03067_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__a22oi_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _00353_ _00355_ _00354_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08123__B1 _00739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10750_ _03471_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07204__B _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4244__B MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09409_ _02021_ _02026_ _02027_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__nand3_2
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10681_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10846__A _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _00299_ _00231_ _00382_ _06537_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__and4_1
XFILLER_205_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08316__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08977__A2 _06604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _05194_ _05195_ _05184_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a21oi_2
XFILLER_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _04064_ _04065_ _04066_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__a21o_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12282_ _05122_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__inv_2
XANTENNA__13183__B1 _04159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11233_ _03991_ _03992_ _03816_ _03862_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a211o_1
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1660_ AuI._0011_ AuI._0012_ AuI._0013_ vssd1 vssd1 vccd1 vccd1 AuI._0014_ sky130_fd_sc_hd__and3_1
XFILLER_106_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _03792_ _03794_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__nand2_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1591_ AuI.pe.Significand\[12\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0765_
+ sky130_fd_sc_hd__or2_1
X_10115_ _02788_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__nor2_2
XFILLER_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11095_ FuI.Integer\[5\] _02931_ _02938_ AuI.result\[5\] _03845_ vssd1 vssd1 vccd1
+ vccd1 _03846_ sky130_fd_sc_hd__a221o_1
XANTENNA__13486__A1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07890__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ _06023_ _02075_ _02020_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__and3b_1
XFILLER_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3550_ MuI._1373_ MuI._1384_ MuI._1395_ vssd1 vssd1 vccd1 vccd1 MuI._1406_ sky130_fd_sc_hd__o21ba_1
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3481_ MuI._0636_ MuI._0394_ MuI._0537_ vssd1 vssd1 vccd1 vccd1 MuI._0647_ sky130_fd_sc_hd__and3_1
XFILLER_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11249__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13116__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11997_ net112 _03593_ _04961_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__and3_1
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5220_ MuI._2860_ MuI._0420_ MuI._0942_ MuI._0941_ vssd1 vssd1 vccd1 vccd1 MuI._0985_
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _03683_ _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__nand2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5151_ MuI._0907_ MuI._0908_ vssd1 vssd1 vccd1 vccd1 MuI._0909_ sky130_fd_sc_hd__nor2_1
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1025_ net107 net33 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0237_ sky130_fd_sc_hd__mux2_1
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _03609_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nand3_1
XMuI._4102_ MuI._2616_ MuI._2850_ vssd1 vssd1 vccd1 vccd1 MuI._3202_ sky130_fd_sc_hd__nand2_1
XMuI._5082_ MuI._2850_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._0833_ sky130_fd_sc_hd__nand2_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08871__D _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ _05482_ _05483_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__o21a_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4033_ MuI._3127_ MuI._3131_ MuI._3132_ vssd1 vssd1 vccd1 vccd1 MuI._3133_ sky130_fd_sc_hd__nand3_1
XFILLER_157_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12549_ _05276_ _05278_ _05277_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__o21bai_1
XFILLER_129_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07640__A2 _04358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__A _02754_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5984_ MuI._1817_ MuI._1825_ vssd1 vssd1 vccd1 vccd1 MuI._1826_ sky130_fd_sc_hd__xnor2_4
XFILLER_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10106__B_N _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4935_ MuI._0666_ MuI._0670_ MuI._0671_ vssd1 vssd1 vccd1 vccd1 MuI._0672_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0809_ AuI._0025_ net114 vssd1 vssd1 vccd1 vccd1 AuI._0029_ sky130_fd_sc_hd__nor2_1
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5512__B1 MuI._3397_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3514__A MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._795_ AuI.pe._399_ AuI.pe._078_ AuI.pe._334_ vssd1 vssd1 vccd1 vccd1 AuI.pe._335_
+ sky130_fd_sc_hd__or3b_1
XFILLER_58_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4866_ MuI._2841_ MuI._3223_ MuI._0478_ MuI._0479_ vssd1 vssd1 vccd1 vccd1 MuI._0596_
+ sky130_fd_sc_hd__o2bb2a_1
X_09760_ _02364_ _02363_ _02355_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a21o_1
XFILLER_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06972_ _05123_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08896__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6605_ MuI._2507_ MuI._2508_ vssd1 vssd1 vccd1 vccd1 MuI._2509_ sky130_fd_sc_hd__nor2_1
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3817_ MuI._2916_ MuI._2704_ MuI._2627_ MuI._2649_ vssd1 vssd1 vccd1 vccd1 MuI._2917_
+ sky130_fd_sc_hd__and4_1
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08711_ _01323_ _01325_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__nand2_1
XMuI._4797_ MuI._0517_ MuI._0518_ MuI._0519_ vssd1 vssd1 vccd1 vccd1 MuI._0520_ sky130_fd_sc_hd__nand3_1
X_09691_ _02147_ _02159_ _02331_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__o211ai_1
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6536_ MuI._2430_ MuI._2431_ vssd1 vssd1 vccd1 vccd1 MuI._2433_ sky130_fd_sc_hd__nor2_1
XFILLER_67_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3748_ MuI._2839_ MuI._2846_ MuI._2842_ vssd1 vssd1 vccd1 vccd1 MuI._2848_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08642_ _01089_ _01088_ _01082_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6467_ MuI._2354_ MuI._2356_ vssd1 vssd1 vccd1 vccd1 MuI._2357_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07305__A net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._3679_ MuI._2517_ MuI._2539_ MuI._2495_ MuI._2550_ vssd1 vssd1 vccd1 vccd1 MuI._2779_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _01187_ _01186_ _01174_ _01135_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__a211oi_1
XANTENNA_MuI._4345__A MuI._0019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5418_ MuI._1188_ MuI._1190_ MuI._1187_ vssd1 vssd1 vccd1 vccd1 MuI._1203_ sky130_fd_sc_hd__o21ba_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07524_ _00121_ _00122_ _00141_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__o21a_1
XMuI._6398_ MuI._2071_ MuI._2280_ vssd1 vssd1 vccd1 vccd1 MuI._2281_ sky130_fd_sc_hd__nor2_1
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5349_ MuI._2895_ MuI._3246_ vssd1 vssd1 vccd1 vccd1 MuI._1127_ sky130_fd_sc_hd__nand2_1
XFILLER_195_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07455_ net50 net51 _04294_ _00072_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__and4_1
XFILLER_211_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10666__A _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12584__C _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08408__A1 _02723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4251__B1 MuI._2352_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _06681_ _00001_ _00003_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__nand3_1
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08136__A _02840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07040__A _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _01740_ _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__or2_1
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11092__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _01672_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__or2_1
XANTENNA__07975__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08007_ _06488_ _05370_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__nand2_1
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10832__C _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07395__A1 _00011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07395__B2 _00012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__A2 _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09958_ _02400_ _02584_ _02620_ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__o211a_1
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08909_ _01521_ _01526_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__xnor2_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07147__A1 _03658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _02491_ _02517_ _02481_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21oi_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _04732_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__nand3_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12121__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_AuI._0943__A0 net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFuI._135__141 vssd1 vssd1 vccd1 vccd1 FuI._135__141/HI net141 sky130_fd_sc_hd__conb_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07215__A _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11851_ _04657_ _04658_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__xor2_1
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _03527_ _03528_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__xnor2_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11782_ _04582_ _04583_ _04572_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a21oi_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _03448_ _03453_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__nand3_1
XFILLER_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13452_ _02921_ _06337_ _02824_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__a21o_1
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10664_ _03222_ _03223_ _03224_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__o21bai_1
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10295__B _02984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ _04994_ _03675_ _02722_ _02916_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__a221o_1
XANTENNA_MuI._5086__A MuI._2919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _06272_ _06273_ _06294_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and3_1
XFILLER_166_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ MuI.result\[2\] _02737_ _02945_ _04004_ _03307_ vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__a221o_1
XFILLER_154_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ _05148_ _05068_ _05177_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand3_1
XANTENNA__07885__A _00502_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ _05093_ _05103_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and3_1
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11706__A1 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11216_ _03970_ _03972_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__and3_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1643_ AuI.exp_a AuI._0710_ AuI._0000_ vssd1 vssd1 vccd1 vccd1 AuI.result\[23\]
+ sky130_fd_sc_hd__a21boi_1
XFILLER_123_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12196_ _02795_ _05028_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or2_1
XANTENNA_MuI._6298__A1 MuI._0801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4720_ MuI._0426_ MuI._0434_ vssd1 vssd1 vccd1 vccd1 MuI._0435_ sky130_fd_sc_hd__xnor2_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 ALU_Output[11] sky130_fd_sc_hd__buf_2
XANTENNA_MuI._6298__B2 MuI._0746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__B _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 ALU_Output[21] sky130_fd_sc_hd__buf_2
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _03898_ _03899_ _03879_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21o_1
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 ALU_Output[31] sky130_fd_sc_hd__buf_2
XAuI._1574_ AuI._0638_ AuI._0749_ vssd1 vssd1 vccd1 vccd1 AuI._0750_ sky130_fd_sc_hd__xnor2_1
XAuI.pe._580_ AuI.pe._125_ AuI.pe._022_ AuI.pe._041_ AuI.pe._105_ AuI.pe._134_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._135_ sky130_fd_sc_hd__a221o_1
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4651_ MuI._0195_ MuI._0358_ vssd1 vssd1 vccd1 vccd1 MuI._0359_ sky130_fd_sc_hd__nand2_1
XANTENNA__09605__A _02377_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11078_ _03513_ _03825_ _03826_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__a21oi_2
XMuI._3602_ MuI._1967_ MuI._1384_ vssd1 vssd1 vccd1 vccd1 MuI._1978_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12131__A1 _00279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3520__A2 MuI._0471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__B2 _00278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4582_ MuI._0014_ MuI._0147_ MuI._0282_ vssd1 vssd1 vccd1 vccd1 MuI._0283_ sky130_fd_sc_hd__nor3_1
X_10029_ _02679_ _02683_ _02697_ _02698_ _02682_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a32o_2
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6321_ MuI._2150_ MuI._2149_ vssd1 vssd1 vccd1 vccd1 MuI._2196_ sky130_fd_sc_hd__or2b_1
XMuI._3533_ MuI._1175_ MuI._1208_ vssd1 vssd1 vccd1 vccd1 MuI._1219_ sky130_fd_sc_hd__or2_1
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11292__D _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6252_ MuI._0361_ MuI._0614_ MuI._3091_ vssd1 vssd1 vccd1 vccd1 MuI._2120_ sky130_fd_sc_hd__and3_1
XFILLER_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3464_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._0460_ sky130_fd_sc_hd__clkbuf_4
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06964__A _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5203_ MuI._0864_ MuI._0858_ MuI._0863_ vssd1 vssd1 vccd1 vccd1 MuI._0967_ sky130_fd_sc_hd__nand3_1
XFILLER_16_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6183_ MuI._2026_ MuI._2027_ MuI._2042_ vssd1 vssd1 vccd1 vccd1 MuI._2045_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6380__A MuI._2789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5134_ MuI._0888_ MuI._0890_ vssd1 vssd1 vccd1 vccd1 MuI._0891_ sky130_fd_sc_hd__nor2_1
X_07240_ _06535_ _06538_ _06536_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o21ai_1
XAuI._1008_ net121 net10 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0220_ sky130_fd_sc_hd__mux2_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5065_ MuI._2841_ MuI._0445_ vssd1 vssd1 vccd1 vccd1 MuI._0815_ sky130_fd_sc_hd__nand2_1
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07171_ _06459_ _06464_ _06462_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__o21ai_1
XFILLER_185_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4016_ MuI._2363_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._3116_ sky130_fd_sc_hd__nand2_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__A _00029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5967_ MuI._1770_ MuI._1793_ MuI._1790_ vssd1 vssd1 vccd1 vccd1 MuI._1807_ sky130_fd_sc_hd__a21o_1
XANTENNA_MuI._4985__D MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4918_ MuI._0613_ MuI._0615_ MuI._0651_ MuI._0652_ vssd1 vssd1 vccd1 vccd1 MuI._0653_
+ sky130_fd_sc_hd__nand4_1
XFILLER_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08122__C _00739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ _02459_ _02460_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a21o_1
XFILLER_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5898_ MuI._1679_ MuI._1720_ MuI._1729_ MuI._1730_ vssd1 vssd1 vccd1 vccd1 MuI._1731_
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._778_ AuI.operand_a\[24\] vssd1 vssd1 vccd1 vccd1 AuI.pe._319_ sky130_fd_sc_hd__inv_2
XFILLER_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4849_ MuI._0574_ MuI._0576_ vssd1 vssd1 vccd1 vccd1 MuI._0577_ sky130_fd_sc_hd__nor2_1
X_06955_ _04940_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[15\] sky130_fd_sc_hd__clkbuf_2
X_09743_ _02380_ _02387_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__nand3_1
XFILLER_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3898__B MuI._2528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _02287_ _02314_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a21boi_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06886_ _04197_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__and3_1
XFILLER_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6519_ MuI._2411_ MuI._2413_ vssd1 vssd1 vccd1 vccd1 MuI._2414_ sky130_fd_sc_hd__nor2_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08625_ _01091_ _01093_ _01104_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__o21a_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12876__A _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08629__A1 _06601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ _01135_ _01136_ _01173_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__nor3_1
XFILLER_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06874__A _04068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__B2 _06606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08792__C _01409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ net51 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__buf_4
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _01091_ _01093_ _01104_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__or3_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _00031_ _00037_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__or2_1
XFILLER_211_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12189__A1 _02862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11004__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07369_ _06662_ _06668_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__and3_1
XFILLER_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ _01373_ _01378_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07604__A2 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _03070_ _03074_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__and3_1
XFILLER_136_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09039_ _01650_ _01651_ _01656_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a21oi_1
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08313__B _00929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__A _00262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__inv_2
XANTENNA_MuI._5353__B MuI._0378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11001_ _02948_ _06562_ _06476_ _00028_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__a22o_1
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _02640_ _05757_ _01962_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a21oi_2
XFILLER_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1290_ AuI._0330_ AuI._0374_ AuI._0263_ vssd1 vssd1 vccd1 vccd1 AuI._0489_ sky130_fd_sc_hd__o21a_1
XANTENNA__12664__A2 _03051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6184__B MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ _04713_ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__xnor2_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _03174_ _05273_ _02745_ _05766_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a311o_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4463__B1 MuI._0019_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ _04640_ _02573_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__xnor2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09817__B1 _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06784__A _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11765_ _04438_ _04439_ _04566_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__a21oi_2
XFILLER_186_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10716_ _03418_ _03435_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__nand3_2
XFILLER_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11696_ _02791_ _04343_ _04492_ _02787_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o211a_1
XFILLER_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13435_ _04011_ _02825_ _06347_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__a211o_1
X_10647_ _03358_ _03361_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__nand3_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13366_ _02820_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xor2_1
XFILLER_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10578_ _03285_ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__xnor2_4
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6870_ MuI._2770_ MuI._2496_ vssd1 vssd1 vccd1 vccd1 MuI._2771_ sky130_fd_sc_hd__xnor2_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12317_ _05159_ _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nor2_1
XFILLER_182_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13297_ _02679_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__or2_2
XFILLER_170_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5821_ MuI._1557_ MuI._1640_ vssd1 vssd1 vccd1 vccd1 MuI._1646_ sky130_fd_sc_hd__nand2_1
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09348__A2 _04509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_AuI.pe._584__A1 AuI.pe._020_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12248_ _05085_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__xor2_4
XFILLER_130_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._701_ AuI.pe._201_ AuI.pe._004_ AuI.pe._040_ AuI.pe._211_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._248_ sky130_fd_sc_hd__a22o_1
XFILLER_170_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5752_ MuI._1500_ MuI._1502_ MuI._1568_ vssd1 vssd1 vccd1 vccd1 MuI._1570_ sky130_fd_sc_hd__nand3_1
XAuI._1626_ AuI._0701_ AuI._0791_ AuI._0792_ AuI._0719_ vssd1 vssd1 vccd1 vccd1 AuI._0793_
+ sky130_fd_sc_hd__a22o_1
X_12179_ FuI.Integer\[13\] _02931_ _03675_ _04865_ _05012_ vssd1 vssd1 vccd1 vccd1
+ _05013_ sky130_fd_sc_hd__a221o_1
XFILLER_122_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI.pe._632_ AuI.pe._074_ AuI.pe._171_ AuI.pe._175_ AuI.pe._183_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe.Significand\[14\] sky130_fd_sc_hd__o22a_1
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06959__A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4703_ MuI._0375_ MuI._0414_ MuI._0415_ vssd1 vssd1 vccd1 vccd1 MuI._0417_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5683_ MuI._1492_ MuI._1493_ vssd1 vssd1 vccd1 vccd1 MuI._1495_ sky130_fd_sc_hd__or2_1
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1557_ AuI._0645_ AuI._0651_ AuI._0663_ AuI._0666_ vssd1 vssd1 vccd1 vccd1 AuI._0736_
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__07781__C _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._563_ AuI.pe._118_ vssd1 vssd1 vccd1 vccd1 AuI.pe._119_ sky130_fd_sc_hd__buf_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4634_ MuI._0335_ MuI._0340_ vssd1 vssd1 vccd1 vccd1 MuI._0341_ sky130_fd_sc_hd__nand2_1
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06740_ _02626_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_49_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1488_ AuI._0537_ AuI._0542_ vssd1 vssd1 vccd1 vccd1 AuI._0674_ sky130_fd_sc_hd__and2_1
XFILLER_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0907__A0 net20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._494_ AuI.pe.significand\[4\] vssd1 vssd1 vccd1 vccd1 AuI.pe._056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4565_ MuI._0077_ MuI._0126_ vssd1 vssd1 vccd1 vccd1 MuI._0265_ sky130_fd_sc_hd__xor2_1
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6304_ MuI._2175_ MuI._2177_ vssd1 vssd1 vccd1 vccd1 MuI._2178_ sky130_fd_sc_hd__xnor2_2
XMuI._3516_ MuI._1021_ vssd1 vssd1 vccd1 vccd1 MuI._1032_ sky130_fd_sc_hd__clkbuf_4
X_08410_ _01022_ _01023_ _01026_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__a21o_1
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4496_ MuI._0055_ MuI._0053_ vssd1 vssd1 vccd1 vccd1 MuI._0189_ sky130_fd_sc_hd__nor2_1
X_09390_ _02004_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__and2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06694__A _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6235_ MuI._2073_ MuI._2074_ MuI._2101_ vssd1 vssd1 vccd1 vccd1 MuI._2102_ sky130_fd_sc_hd__nand3_1
XANTENNA__09070__A _06488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3447_ MuI._0229_ MuI._0251_ MuI._0262_ vssd1 vssd1 vccd1 vccd1 MuI._0273_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _06463_ _05305_ _05370_ _06492_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__a22oi_2
XANTENNA__11615__B1 _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4623__A MuI.b_operand\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6166_ MuI._2018_ MuI._2024_ MuI._2025_ vssd1 vssd1 vccd1 vccd1 MuI._2026_ sky130_fd_sc_hd__nand3_1
X_08272_ _00575_ _00576_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11091__B2 _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._3884__D MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5117_ MuI._0848_ MuI._0850_ MuI._0849_ vssd1 vssd1 vccd1 vccd1 MuI._0872_ sky130_fd_sc_hd__o21bai_1
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._710__A AuI.pe.significand\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07223_ _06499_ _06502_ _06505_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__o21ba_1
XANTENNA__08117__C _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6097_ MuI._0625_ MuI._2797_ MuI._2789_ MuI._0372_ vssd1 vssd1 vccd1 vccd1 MuI._1950_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5048_ MuI.a_operand\[8\] MuI.a_operand\[7\] MuI._2884_ MuI._2880_ vssd1 vssd1
+ vccd1 vccd1 MuI._0796_ sky130_fd_sc_hd__and4_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _06453_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__xnor2_2
XFILLER_180_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5706__B1 MuI._3185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ _04736_ _06284_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__and2_1
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07675__D _06443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5173__B MuI._2854_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12343__A1 _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11775__A _00345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 net53 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_4
Xfanout124 net32 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_4
XFILLER_160_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06869__A _04015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input1_A Operation[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08787__C _03960_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07987_ _00299_ _00231_ _06433_ _00287_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__and4_1
XANTENNA__07691__C net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5485__A2 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3702__A MuI._2693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09726_ _02431_ _02229_ net115 _06436_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__and4_1
X_06938_ net9 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__buf_2
XFILLER_68_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4517__B MuI._2918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06869_ _04015_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[1\] sky130_fd_sc_hd__buf_2
X_09657_ _06463_ _00592_ _00072_ _06492_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22oi_2
XANTENNA_AuI._0933__A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08608_ _01218_ _01224_ _01225_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__a21o_1
X_09588_ _06560_ _06443_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__nand2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4996__A1 MuI._0636_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__D _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13214__B _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08539_ _01143_ _01142_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__and2_1
XFILLER_169_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08078__A2 _00259_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08308__B _00919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11550_ _04161_ _04328_ _04333_ _04335_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__a211o_1
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07825__A2 _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _03203_ _03204_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a21o_1
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6170__D MuI._2803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _04259_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__xor2_2
XFILLER_149_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ _06125_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__and2_1
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ _02020_ _06023_ _02140_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and3_1
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13151_ _06015_ _05971_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _00756_ _00758_ _00757_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__o21bai_1
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _04793_ _04795_ _04794_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__o21bai_1
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _05979_ _05980_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input57_A b_operand[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _03432_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__buf_4
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08978__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _04815_ _04853_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__and3_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12885__A2 _05758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06779__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0827__B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1411_ AuI._0597_ AuI._0598_ AuI._0599_ vssd1 vssd1 vccd1 vccd1 AuI.pe.significand\[24\]
+ sky130_fd_sc_hd__a21oi_4
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3612__A MuI._2077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1342_ AuI._0389_ AuI._0295_ AuI._0422_ vssd1 vssd1 vccd1 vccd1 AuI._0537_ sky130_fd_sc_hd__and3_1
XFILLER_92_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13295__C1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4427__B MuI._0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__C _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A2 _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12935_ _05822_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nor2_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1273_ AuI._0389_ AuI._0471_ AuI._0421_ AuI._0472_ vssd1 vssd1 vccd1 vccd1 AuI._0473_
+ sky130_fd_sc_hd__o211a_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4350_ MuI._1032_ MuI._2886_ MuI._2882_ MuI._0790_ vssd1 vssd1 vccd1 vccd1 MuI._0029_
+ sky130_fd_sc_hd__a22oi_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ _05565_ _05665_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__nor2_1
XFILLER_206_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI._0893__B_N net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4281_ MuI._2822_ MuI._3235_ MuI._3240_ MuI._3250_ vssd1 vssd1 vccd1 vccd1 MuI._3381_
+ sky130_fd_sc_hd__o31a_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _02790_ _04349_ _01350_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__o21a_1
XFILLER_187_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6020_ MuI._0735_ MuI._1153_ MuI._2682_ MuI._2594_ vssd1 vssd1 vccd1 vccd1 MuI._1865_
+ sky130_fd_sc_hd__and4_1
XFILLER_159_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12797_ _05209_ _02941_ _02731_ AuI.result\[19\] vssd1 vssd1 vccd1 vccd1 _05677_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07122__B _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _04398_ _04419_ _04547_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a211oi_2
XFILLER_159_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI.pe._530__A AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10764__A _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11679_ _04250_ _04364_ _04473_ _04474_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__a211oi_4
XFILLER_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13418_ _06330_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__nand2_1
XFILLER_162_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08234__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _02683_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__xor2_4
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0988_ AuI._0168_ vssd1 vssd1 vccd1 vccd1 AuI._0200_ sky130_fd_sc_hd__clkbuf_2
XFILLER_170_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6853_ MuI._2758_ vssd1 vssd1 vccd1 vccd1 MuI.result\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._557__B2 AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5804_ MuI._1624_ MuI._1625_ MuI._1536_ MuI._1597_ vssd1 vssd1 vccd1 vccd1 MuI._1628_
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6784_ MuI._2568_ MuI._2571_ MuI._2575_ vssd1 vssd1 vccd1 vccd1 MuI._2706_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07910_ _00524_ _00526_ _00525_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a21o_1
XMuI._3996_ MuI._3093_ MuI._3094_ MuI._3095_ vssd1 vssd1 vccd1 vccd1 MuI._3096_ sky130_fd_sc_hd__nand3b_1
X_08890_ _01470_ _01481_ _01506_ _01507_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a211oi_2
XANTENNA__06689__A _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5735_ MuI._0990_ MuI._1550_ MuI._1551_ vssd1 vssd1 vccd1 vccd1 MuI._1552_ sky130_fd_sc_hd__and3_1
XFILLER_97_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1609_ AuI._0670_ AuI._0673_ vssd1 vssd1 vccd1 vccd1 AuI._0779_ sky130_fd_sc_hd__or2b_1
XANTENNA__07201__B1 _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07841_ _03324_ _04456_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__nand2_1
XAuI.pe._615_ AuI.pe._145_ AuI.pe._141_ AuI.pe._158_ vssd1 vssd1 vccd1 vccd1 AuI.pe._168_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_AuI.pe._408__C AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5666_ MuI._1009_ MuI._1466_ MuI._1475_ vssd1 vssd1 vccd1 vccd1 MuI._1476_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._3522__A MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _00159_ _00167_ _00158_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a21bo_1
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._546_ AuI.pe._101_ AuI.pe._103_ AuI.pe._074_ vssd1 vssd1 vccd1 vccd1 AuI.pe._104_
+ sky130_fd_sc_hd__a21o_1
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4617_ MuI._0321_ MuI._0449_ vssd1 vssd1 vccd1 vccd1 MuI._0322_ sky130_fd_sc_hd__nand2_1
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06723_ _02442_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__and3_1
X_09511_ _02120_ _02123_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a211oi_1
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5597_ MuI._1393_ MuI._1397_ MuI._1398_ MuI._1399_ vssd1 vssd1 vccd1 vccd1 MuI._1400_
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._477_ AuI.pe._040_ vssd1 vssd1 vccd1 vccd1 AuI.pe._041_ sky130_fd_sc_hd__buf_2
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4548_ MuI._0245_ vssd1 vssd1 vccd1 vccd1 MuI._0246_ sky130_fd_sc_hd__buf_4
X_09442_ _06579_ net127 _06431_ _06578_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a22oi_2
XFILLER_37_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4978__A1 MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4479_ MuI._2605_ MuI._2873_ MuI._2875_ MuI._2852_ vssd1 vssd1 vccd1 vccd1 MuI._0170_
+ sky130_fd_sc_hd__a22oi_1
X_09373_ _01965_ _01980_ _01979_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a21o_1
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6218_ MuI._2041_ MuI._2075_ MuI._2082_ vssd1 vssd1 vccd1 vccd1 MuI._2083_ sky130_fd_sc_hd__and3_1
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10377__C _00382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ _00939_ _00940_ _00933_ _00936_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__o211ai_2
XFILLER_178_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4072__B MuI._3171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6149_ MuI._0504_ MuI._2006_ vssd1 vssd1 vccd1 vccd1 MuI._2007_ sky130_fd_sc_hd__and2_1
XFILLER_165_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10811__A1 _03443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _00641_ _00642_ _00561_ _00643_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__or4bb_2
XANTENNA__10811__B2 _00281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07206_ _06499_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _00749_ _00803_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__xor2_2
XANTENNA__07686__C _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ _06432_ _06435_ net58 _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__and4bb_1
XFILLER_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07983__A _00313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _04197_ _06067_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__and2_1
XANTENNA__13108__A3 _06000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11119__A2 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10613__S _02926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13209__B _05713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._6373__A1_N MuI._0867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12619__A2 _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _02350_ _02351_ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a21bo_1
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10981_ _03716_ _03719_ _03720_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__nand3_2
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10849__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ _05134_ _03067_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__and2b_1
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09422__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ _05517_ _05518_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xor2_1
XFILLER_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4263__A MuI._3362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _04386_ _04389_ _04390_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__nand3_1
XANTENNA__11055__A1 _02485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5078__B MuI._2838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12582_ _05270_ _05274_ _05271_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__o21bai_1
XANTENNA__11055__B2 _06565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ _04150_ _04152_ _04023_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__o21a_1
XFILLER_156_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._157_ FuI.a_operand\[27\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[27\] sky130_fd_sc_hd__clkbuf_1
XAuI._0911_ net113 AuI._0128_ AuI._0129_ vssd1 vssd1 vccd1 vccd1 AuI._0130_ sky130_fd_sc_hd__and3_1
X_11464_ _04041_ _04043_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__nand2_1
XFILLER_184_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._088_ FuI.a_operand\[6\] FuI._050_ vssd1 vssd1 vccd1 vccd1 FuI._051_ sky130_fd_sc_hd__and2_1
X_10415_ _00807_ _00808_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__nand2_1
X_13203_ _06017_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__o21ba_1
XAuI._0842_ net126 vssd1 vssd1 vccd1 vccd1 AuI._0062_ sky130_fd_sc_hd__inv_2
X_11395_ MuI.result\[7\] _02737_ _02945_ _04327_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__08223__A2 _06584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ _03006_ _00768_ _03038_ _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211o_1
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ _03507_ _05906_ _05981_ _03454_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__a22oi_1
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0838__A net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3850_ MuI._2945_ MuI._2948_ vssd1 vssd1 vccd1 vccd1 MuI._2950_ sky130_fd_sc_hd__nor2_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13065_ _05961_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__and2_1
XFILLER_79_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10318__B1 _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ net58 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__clkbuf_4
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _00292_ _00534_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a22o_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3781_ MuI._2880_ vssd1 vssd1 vccd1 vccd1 MuI._2881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5520_ MuI._2876_ MuI._0245_ MuI._0320_ MuI._2874_ vssd1 vssd1 vccd1 vccd1 MuI._1315_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._400_ AuI.pe.significand\[16\] vssd1 vssd1 vccd1 vccd1 AuI.pe._367_ sky130_fd_sc_hd__buf_2
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5451_ MuI._1181_ MuI._1238_ vssd1 vssd1 vccd1 vccd1 MuI._1239_ sky130_fd_sc_hd__nor2_1
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._525__A AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1325_ AuI._0520_ AuI._0521_ vssd1 vssd1 vccd1 vccd1 AuI._0522_ sky130_fd_sc_hd__nor2_2
XFILLER_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09487__A1 _06548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4402_ MuI.a_operand\[7\] vssd1 vssd1 vccd1 vccd1 MuI._0085_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09487__B2 _02291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5382_ MuI._1161_ MuI._1162_ vssd1 vssd1 vccd1 vccd1 MuI._1163_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12918_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__nor2_1
XAuI._1256_ AuI._0435_ AuI._0445_ AuI._0446_ vssd1 vssd1 vccd1 vccd1 AuI._0458_ sky130_fd_sc_hd__o21a_1
XANTENNA_MuI._3880__A1 MuI._2066_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4333_ MuI._0006_ MuI._0008_ vssd1 vssd1 vccd1 vccd1 MuI._0011_ sky130_fd_sc_hd__nor2_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07133__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13035__A2 _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1187_ AuI._0367_ AuI._0382_ AuI._0392_ vssd1 vssd1 vccd1 vccd1 AuI._0393_ sky130_fd_sc_hd__a21o_1
X_12849_ _05629_ _05646_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__nor2_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4264_ MuI._1142_ MuI._2374_ MuI._3363_ MuI._2939_ vssd1 vssd1 vccd1 vccd1 MuI._3364_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06972__A _05123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6003_ MuI._1843_ MuI._1845_ vssd1 vssd1 vccd1 vccd1 MuI._1847_ sky130_fd_sc_hd__xor2_2
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4195_ MuI._3176_ MuI._3177_ vssd1 vssd1 vccd1 vccd1 MuI._3295_ sky130_fd_sc_hd__xor2_1
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12185__S _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__A _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08462__A2 _00074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08040_ _00255_ _00256_ _00368_ _00369_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__and4_1
XFILLER_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11349__A2 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3517__A MuI._1032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10644__D _00059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09991_ _01311_ _01312_ _01313_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__or3_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6836_ MuI._2750_ vssd1 vssd1 vccd1 vccd1 MuI.result\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_130_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ _01551_ _01552_ _01559_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a21o_1
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07953__D _00047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__B _04531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6767_ MuI._2685_ MuI._2596_ MuI._2600_ MuI._2686_ vssd1 vssd1 vccd1 vccd1 MuI._2687_
+ sky130_fd_sc_hd__or4_1
XFILLER_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3979_ MuI._2994_ MuI._3077_ MuI._3078_ vssd1 vssd1 vccd1 vccd1 MuI._3079_ sky130_fd_sc_hd__or3_1
XFILLER_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08873_ _01487_ _01490_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__xnor2_1
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1223__C1 AuI._0139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5718_ MuI._1530_ MuI._1531_ MuI._1525_ vssd1 vssd1 vccd1 vccd1 MuI._1533_ sky130_fd_sc_hd__a21o_1
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6698_ MuI._0999_ MuI._2482_ MuI._2483_ MuI._2607_ vssd1 vssd1 vccd1 vccd1 MuI._2611_
+ sky130_fd_sc_hd__o31a_1
X_07824_ _00219_ _00220_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__nand2_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5649_ MuI._1242_ MuI._1331_ MuI._1454_ MuI._1456_ vssd1 vssd1 vccd1 vccd1 MuI._1457_
+ sky130_fd_sc_hd__o22a_1
XFILLER_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07755_ _00168_ _00169_ _00170_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__and3_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._529_ AuI.pe._046_ AuI.pe._054_ AuI.pe._087_ vssd1 vssd1 vccd1 vccd1 AuI.pe._088_
+ sky130_fd_sc_hd__a21o_1
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06706_ _02259_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__and3_1
X_07686_ _00300_ _00302_ _00270_ _00303_ vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__and4bb_1
XANTENNA__08139__A _06578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__A _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5179__A MuI._2583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09425_ _02043_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__nor2_1
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5612__A2 MuI._0112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI.pe._466__B1 AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _06495_ net7 _00032_ _06494_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a22oi_2
XANTENNA__06882__A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _00596_ _00919_ _00924_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__a21o_1
X_09287_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08238_ _00852_ _00855_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__or2b_1
XFILLER_193_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._769__A1 AuI.pe._056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12537__A1 _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ _00784_ _00786_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__nor2_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _02715_ _02753_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a21bo_1
XFILLER_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11180_ _03934_ _03935_ _03926_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__a21o_1
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08602__A net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11760__A2 _04725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _05338_ _03239_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__or2b_1
XFILLER_122_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10062_ _04004_ _02719_ _02725_ _02733_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a211o_1
XANTENNA__07218__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12882__A1_N _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5080__C MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07192__A2 _06466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09433__A _06520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__A1 _02205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09469__B2 _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1110_ AuI._0319_ vssd1 vssd1 vccd1 vccd1 AuI._0320_ sky130_fd_sc_hd__clkbuf_2
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09152__B _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ _03525_ _04380_ _03522_ _03521_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__a31o_2
XANTENNA__10298__B _04380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ _05575_ _05572_ _02607_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__a21o_1
XAuI._1041_ AuI._0140_ AuI._0252_ vssd1 vssd1 vccd1 vccd1 AuI._0253_ sky130_fd_sc_hd__nand2_1
XANTENNA__10729__D _05820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ _03621_ _03628_ _03629_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nand3_1
XFILLER_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07888__A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12634_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and2b_1
XANTENNA__06792__A _03174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0840__B net116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4143__D MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ _05425_ _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__nor2_1
XFILLER_157_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._5367__A1 MuI._2869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__A_N _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5367__B2 MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _04296_ _04297_ _04094_ _04183_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o211a_1
XFILLER_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ _04999_ _04996_ _05353_ _05350_ _05351_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__o2111a_1
XANTENNA_MuI._4440__B MuI._0076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _02658_ _03082_ _00789_ _06585_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__a22o_1
XFILLER_153_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4951_ MuI._0686_ MuI._0688_ vssd1 vssd1 vccd1 vccd1 MuI._0689_ sky130_fd_sc_hd__or2b_1
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0825_ AuI._0036_ net13 AuI._0044_ net133 vssd1 vssd1 vccd1 vccd1 AuI._0045_
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _03997_ _03999_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nor2_2
XANTENNA_output88_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3902_ MuI._2998_ MuI._2999_ MuI._3001_ vssd1 vssd1 vccd1 vccd1 MuI._3002_ sky130_fd_sc_hd__nand3b_1
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07955__A1 _00062_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07955__B2 _00063_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5552__A MuI._3268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4882_ MuI._0588_ MuI._0611_ MuI._0612_ MuI._0528_ vssd1 vssd1 vccd1 vccd1 MuI._0613_
+ sky130_fd_sc_hd__a211o_1
X_10329_ _00727_ _00059_ _04714_ _00728_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a22oi_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _06016_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6621_ MuI._1446_ MuI._1430_ vssd1 vssd1 vccd1 vccd1 MuI._2526_ sky130_fd_sc_hd__or2b_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3833_ MuI._2929_ MuI._2932_ vssd1 vssd1 vccd1 vccd1 MuI._2933_ sky130_fd_sc_hd__xor2_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07128__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _03497_ _05831_ _05941_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and4_1
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6552_ MuI._2185_ MuI._2204_ vssd1 vssd1 vccd1 vccd1 MuI._2450_ sky130_fd_sc_hd__or2_1
XANTENNA__12161__C1 _04992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3764_ MuI._2858_ MuI._2859_ MuI._2863_ vssd1 vssd1 vccd1 vccd1 MuI._2864_ sky130_fd_sc_hd__nand3_1
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5503_ MuI._1258_ MuI._1257_ MuI._1249_ vssd1 vssd1 vccd1 vccd1 MuI._1297_ sky130_fd_sc_hd__a21o_1
XANTENNA__06967__A _05058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6483_ MuI._1919_ MuI._1920_ MuI._2373_ vssd1 vssd1 vccd1 vccd1 MuI._2375_ sky130_fd_sc_hd__o21ai_2
XFILLER_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3695_ MuI._2759_ MuI._2779_ MuI._2778_ vssd1 vssd1 vccd1 vccd1 MuI._2795_ sky130_fd_sc_hd__o21ai_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5434_ MuI._2976_ MuI._0246_ MuI._0321_ MuI._2975_ vssd1 vssd1 vccd1 vccd1 MuI._1221_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3800__A MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._6814__C MuI._2733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _00155_ _00156_ _00157_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__nand3_1
XAuI._1308_ net10 net42 AuI._0125_ vssd1 vssd1 vccd1 vccd1 AuI._0506_ sky130_fd_sc_hd__mux2_2
XFILLER_207_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5365_ MuI._1140_ MuI._1144_ vssd1 vssd1 vccd1 vccd1 MuI._1145_ sky130_fd_sc_hd__xnor2_1
XAuI._1239_ AuI._0425_ AuI._0440_ vssd1 vssd1 vccd1 vccd1 AuI._0442_ sky130_fd_sc_hd__and2_1
X_07471_ net34 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__buf_4
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4316_ MuI._3413_ MuI._3415_ vssd1 vssd1 vccd1 vccd1 MuI._3416_ sky130_fd_sc_hd__xor2_2
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _01825_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nand3_1
XFILLER_210_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5296_ MuI._0085_ MuI._3306_ MuI.a_operand\[6\] MuI._3307_ vssd1 vssd1 vccd1
+ vccd1 MuI._1069_ sky130_fd_sc_hd__and4_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4247_ MuI._3346_ MuI._3226_ vssd1 vssd1 vccd1 vccd1 MuI._3347_ sky130_fd_sc_hd__xnor2_1
X_09141_ _01415_ _01435_ _01434_ _01431_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__o211a_1
XANTENNA__12209__A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11113__A _03713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4178_ MuI._3257_ MuI._3276_ MuI._3277_ vssd1 vssd1 vccd1 vccd1 MuI._3278_ sky130_fd_sc_hd__a21oi_2
X_09072_ _06494_ _00150_ net10 net11 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__and4_1
XFILLER_175_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12519__A1 _03134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08023_ _00635_ _00638_ _00639_ _00640_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a211oi_4
XANTENNA_MuI._4030__A1 MuI._0570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4030__B2 MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11767__B _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08779__D _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _01767_ _01959_ _01963_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__and3_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6819_ MuI._2740_ vssd1 vssd1 vccd1 vccd1 MuI.result\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07038__A _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _01540_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08856_ _06663_ _00048_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nand2_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__A _01203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07807_ _06606_ _06601_ _05112_ _05187_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__and4_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4228__D MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08787_ _00921_ _01206_ _03960_ _06446_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__and4_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ _00353_ _00354_ _00355_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__and3_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07204__C _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07669_ _04165_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__clkbuf_4
X_09408_ _02019_ _02018_ _02017_ _01995_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a211o_1
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10680_ _03324_ _04714_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nand2_1
XANTENNA__13404__C1 _02750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10846__B _04789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ _01952_ _01955_ _01925_ _01840_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a211oi_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__B _03928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _05184_ _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__and3_2
XFILLER_193_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _04064_ _04065_ _04066_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand3_2
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12281_ _05035_ _04981_ _05120_ _05121_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__a211oi_4
XFILLER_107_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13183__A1 _02645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ _03816_ _03862_ _03991_ _03992_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o211a_1
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11163_ _03916_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nor2_1
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1590_ AuI._0693_ AuI._0757_ AuI._0763_ AuI._0703_ vssd1 vssd1 vccd1 vccd1 AuI._0764_
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10114_ _02604_ _04542_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and2b_1
XFILLER_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ MuI.result\[5\] _02737_ _02945_ _04197_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13486__A2 _06394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _02708_ _02711_ _02713_ _02714_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a32o_1
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13238__A2 _06045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3480_ MuI._0625_ vssd1 vssd1 vccd1 vccd1 MuI._0636_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11249__A1 _02129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11996_ _04510_ _04694_ _04695_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__nand3_1
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ _02769_ _03321_ _03684_ _03317_ _02762_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__a2111o_1
XFILLER_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0851__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5150_ MuI._0477_ MuI._2765_ MuI._3306_ MuI._3307_ vssd1 vssd1 vccd1 vccd1 MuI._0908_
+ sky130_fd_sc_hd__and4_1
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1024_ AuI._0192_ vssd1 vssd1 vccd1 vccd1 AuI._0236_ sky130_fd_sc_hd__buf_2
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4101_ MuI._3198_ MuI._3199_ MuI._3200_ vssd1 vssd1 vccd1 vccd1 MuI._3201_ sky130_fd_sc_hd__o21ba_1
X_10878_ _03428_ _03426_ _03427_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__a21bo_1
XFILLER_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5081_ MuI._0829_ MuI._0831_ vssd1 vssd1 vccd1 vccd1 MuI._0832_ sky130_fd_sc_hd__nor2_1
XANTENNA__07411__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _05482_ _05483_ _06427_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__a21oi_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12029__A _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4032_ MuI._3129_ MuI._3130_ MuI._3128_ vssd1 vssd1 vccd1 vccd1 MuI._3132_ sky130_fd_sc_hd__a21bo_1
XFILLER_200_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ _00262_ _03257_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a22o_1
XFILLER_157_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__A _00125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _05226_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or3_4
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5983_ MuI._1818_ MuI._1822_ MuI._1823_ vssd1 vssd1 vccd1 vccd1 MuI._1825_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11587__B _02797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6378__A MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4934_ MuI._0502_ MuI._0544_ vssd1 vssd1 vccd1 vccd1 MuI._0671_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0808_ net50 AuI._0026_ net49 AuI._0027_ vssd1 vssd1 vccd1 vccd1 AuI._0028_ sky130_fd_sc_hd__o22a_1
XANTENNA_MuI._5713__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI.pe._794_ AuI.pe.significand\[20\] AuI.pe._368_ AuI.pe._076_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._334_ sky130_fd_sc_hd__or3_1
XFILLER_101_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4865_ MuI._0591_ MuI._0594_ vssd1 vssd1 vccd1 vccd1 MuI._0595_ sky130_fd_sc_hd__nor2_1
XFILLER_140_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06971_ _05112_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__buf_4
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3816_ MuI._2840_ vssd1 vssd1 vccd1 vccd1 MuI._2916_ sky130_fd_sc_hd__buf_2
XMuI._6604_ MuI._1839_ MuI._1836_ vssd1 vssd1 vccd1 vccd1 MuI._2508_ sky130_fd_sc_hd__and2b_1
XANTENNA__08896__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _00951_ _00953_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__xnor2_2
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4796_ MuI._0469_ MuI._0472_ vssd1 vssd1 vccd1 vccd1 MuI._0519_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09690_ _01996_ _02014_ _02015_ _02016_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__nand4_1
XANTENNA__06697__A _02118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6535_ MuI._2430_ MuI._2431_ vssd1 vssd1 vccd1 vccd1 MuI._2432_ sky130_fd_sc_hd__and2_1
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3747_ MuI._2839_ MuI._2842_ MuI._2846_ vssd1 vssd1 vccd1 vccd1 MuI._2847_ sky130_fd_sc_hd__or3_1
XFILLER_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08641_ _01089_ _01082_ _01088_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__and3_1
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._669__B1 AuI.pe._023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6466_ MuI._2318_ MuI._2355_ vssd1 vssd1 vccd1 vccd1 MuI._2356_ sky130_fd_sc_hd__nand2_1
XMuI._3678_ MuI._1263_ MuI._2773_ vssd1 vssd1 vccd1 vccd1 MuI._2778_ sky130_fd_sc_hd__nand2_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ _01137_ _01155_ _01189_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__o21a_1
XFILLER_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5417_ MuI._1184_ MuI._1185_ MuI._1201_ vssd1 vssd1 vccd1 vccd1 MuI._1202_ sky130_fd_sc_hd__nand3_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6397_ MuI._2067_ MuI._2070_ vssd1 vssd1 vccd1 vccd1 MuI._2280_ sky130_fd_sc_hd__nor2_1
X_07523_ _00129_ _00140_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__xnor2_4
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5348_ MuI._1124_ MuI._1125_ vssd1 vssd1 vccd1 vccd1 MuI._1126_ sky130_fd_sc_hd__nor2_1
XFILLER_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13323__A _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07454_ net34 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__buf_4
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10666__B _00216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5457__A MuI._3306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5279_ MuI._1029_ MuI._1048_ MuI._1049_ vssd1 vssd1 vccd1 vccd1 MuI._1050_ sky130_fd_sc_hd__and3_1
XANTENNA__12584__D _03424_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07385_ _00000_ _06682_ _00002_ _06568_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nand4_1
XANTENNA_MuI._4251__B2 MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08408__A2 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__B _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09124_ _01426_ _01741_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nor2_2
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _01665_ _01666_ _01671_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__o21ba_1
XFILLER_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07975__B net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09369__B1 _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08006_ _06496_ _06493_ _06490_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__o21ai_1
XFILLER_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10832__D _00412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07395__A2 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _02324_ _02346_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__nand2_1
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _01524_ _01525_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__nor2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _02524_ _02518_ _02525_ _02545_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__or4_2
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07147__A2 _03873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _06460_ _06604_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__and2_1
XFILLER_206_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4536__A MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__B _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0943__A1 net23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11850_ _02862_ _05831_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nand2_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ _03722_ _04316_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__and2_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04572_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__and3_1
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07855__B1 _00471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _03452_ _03451_ _03450_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13451_ _06364_ _06170_ _06342_ _06365_ _02711_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__a311o_1
XFILLER_9_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ _03221_ _03236_ _03237_ _03241_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__a31o_1
XANTENNA__10295__C _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _02916_ _04929_ _02744_ _04627_ FuI.Integer\[15\] vssd1 vssd1 vccd1 vccd1
+ _05253_ sky130_fd_sc_hd__a32o_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._5086__B MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ _04068_ _02727_ _02767_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__o22ai_1
X_13382_ _06272_ _06273_ _06294_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__a21oi_1
XFILLER_194_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ _05148_ _05068_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a21o_1
XANTENNA__07885__B _03917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09158__A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12264_ _05102_ _05099_ _05100_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__nand3_2
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10205__A_N _02442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1642_ AuI.exponent_sub\[0\] AuI._0769_ AuI._0708_ AuI.exp_a AuI._0699_ vssd1
+ vssd1 vccd1 vccd1 AuI._0000_ sky130_fd_sc_hd__o221a_1
X_11215_ _03163_ _00421_ _03762_ _03973_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a32o_1
X_12195_ _02795_ _05028_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__nand2_1
XFILLER_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._6298__A2 MuI._1164_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__C _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 ALU_Output[12] sky130_fd_sc_hd__buf_2
XFILLER_150_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1573_ AuI._0639_ AuI._0745_ AuI._0641_ vssd1 vssd1 vccd1 vccd1 AuI._0749_ sky130_fd_sc_hd__a21oi_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 ALU_Output[22] sky130_fd_sc_hd__buf_2
X_11146_ _03879_ _03898_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nand3_1
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 ALU_Output[3] sky130_fd_sc_hd__buf_2
XFILLER_150_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4650_ MuI._0192_ MuI._0194_ vssd1 vssd1 vccd1 vccd1 MuI._0358_ sky130_fd_sc_hd__or2_1
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09605__B _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11077_ _03647_ _03649_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__nor2_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3601_ MuI._1395_ MuI._1373_ vssd1 vssd1 vccd1 vccd1 MuI._1967_ sky130_fd_sc_hd__nor2_1
XFILLER_209_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12131__A2 _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4581_ MuI._0148_ MuI._0281_ vssd1 vssd1 vccd1 vccd1 MuI._0282_ sky130_fd_sc_hd__xnor2_1
X_10028_ _02665_ _02677_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__nand2_1
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6320_ MuI._2193_ MuI._2155_ vssd1 vssd1 vccd1 vccd1 MuI._2195_ sky130_fd_sc_hd__xor2_1
XFILLER_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3532_ MuI._0592_ MuI._0889_ MuI._1197_ vssd1 vssd1 vccd1 vccd1 MuI._1208_ sky130_fd_sc_hd__and3_1
XFILLER_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12419__B1 _03449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6251_ MuI._2117_ MuI._2118_ vssd1 vssd1 vccd1 vccd1 MuI._2119_ sky130_fd_sc_hd__nor2_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3463_ MuI._0438_ vssd1 vssd1 vccd1 vccd1 MuI._0449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._520__C1 AuI.pe._037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5202_ MuI._0961_ MuI._0963_ MuI._0964_ vssd1 vssd1 vccd1 vccd1 MuI._0965_ sky130_fd_sc_hd__a21bo_1
X_11979_ _04793_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__o21ai_1
XFILLER_189_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6182_ MuI._2026_ MuI._2027_ MuI._2042_ vssd1 vssd1 vccd1 vccd1 MuI._2043_ sky130_fd_sc_hd__and3_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5133_ MuI._2869_ MuI._0088_ MuI._2319_ MuI._2867_ vssd1 vssd1 vccd1 vccd1 MuI._0890_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_MuI._6380__B MuI._0438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI._1007_ AuI._0190_ AuI._0191_ AuI._0218_ vssd1 vssd1 vccd1 vccd1 AuI._0219_ sky130_fd_sc_hd__or3b_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4181__A MuI._3278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5064_ MuI._0811_ MuI._0813_ vssd1 vssd1 vccd1 vccd1 MuI._0814_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._4612__C MuI._0315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07170_ _06467_ _06468_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__o21bai_1
XFILLER_158_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06980__A _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4015_ MuI._3113_ MuI._3114_ vssd1 vssd1 vccd1 vccd1 MuI._3115_ sky130_fd_sc_hd__nor2_1
XFILLER_200_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__B _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5966_ MuI._1804_ MuI._1805_ vssd1 vssd1 vccd1 vccd1 MuI._1806_ sky130_fd_sc_hd__nor2_1
XFILLER_160_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4917_ MuI._0649_ MuI._0650_ MuI._0633_ MuI._0646_ vssd1 vssd1 vccd1 vccd1 MuI._0652_
+ sky130_fd_sc_hd__a211o_1
X_09811_ _02248_ _04035_ _02461_ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a31o_1
XMuI._5897_ MuI._1724_ MuI._1726_ MuI._1728_ MuI._0727_ vssd1 vssd1 vccd1 vccd1 MuI._1730_
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._777_ AuI.pe._377_ AuI.pe._381_ AuI.pe._398_ AuI.pe._018_ AuI.exp_a vssd1
+ vssd1 vccd1 vccd1 AuI.pe._318_ sky130_fd_sc_hd__a41o_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4848_ MuI._0574_ MuI._0575_ MuI._2484_ MuI.b_operand\[8\] vssd1 vssd1 vccd1
+ vccd1 MuI._0576_ sky130_fd_sc_hd__and4bb_1
X_09742_ _02385_ _02386_ _02376_ _02384_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a211o_1
X_06954_ _04929_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__and3_1
XANTENNA__12222__A _00921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4779_ MuI._0497_ MuI._0499_ vssd1 vssd1 vccd1 vccd1 MuI._0500_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09673_ _02309_ _02312_ _02263_ _02288_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__o211ai_1
X_06885_ _04186_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__buf_4
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6518_ MuI._2143_ MuI._2412_ vssd1 vssd1 vccd1 vccd1 MuI._2413_ sky130_fd_sc_hd__or2_1
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _01236_ _01240_ _01228_ _01241_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__o211ai_4
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12876__B _05209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._443__A AuI.pe.significand\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6449_ MuI._2309_ MuI._2331_ MuI._2336_ vssd1 vssd1 vccd1 vccd1 MuI._2337_ sky130_fd_sc_hd__nor3_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _01156_ _01172_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08629__A2 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07506_ net50 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__buf_4
XFILLER_211_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08486_ _01096_ _01103_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07051__A _05970_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07437_ _00052_ _00054_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__nand2_1
XFILLER_196_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4091__A MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12189__A2 _04865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ _06665_ _06667_ _06664_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06890__A _04240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _01705_ _01701_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__or2b_1
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07299_ _06598_ _06599_ _04832_ _04896_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__and4_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09038_ _01653_ _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__xnor2_1
XFILLER_164_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11020__B _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12897__B1 _05981_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _03600_ _03603_ _03601_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09706__A _06504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09762__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12132__A _03378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07226__A _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _05838_ _05839_ _03133_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__o21a_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11971__A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ _03722_ _04800_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__and2_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _05273_ _02727_ _02738_ MuI.result\[20\] vssd1 vssd1 vccd1 vccd1 _05768_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _02574_ _02521_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2b_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5660__B1 MuI._0420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4942__A2_N MuI._0168_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__B1 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__B1 _05700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04436_ _04437_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__and2_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10715_ _03433_ _03434_ _03423_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__a21o_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _02789_ _02785_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__or2b_1
XFILLER_186_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13434_ MuI.result\[29\] _02736_ _02730_ AuI.result\[29\] _06348_ vssd1 vssd1 vccd1
+ vccd1 _06349_ sky130_fd_sc_hd__a221o_1
XFILLER_139_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10646_ _02987_ _04531_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__nand4_1
X_13365_ _03680_ _05992_ _06108_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__and3_1
X_10577_ _02954_ _03286_ _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a21oi_2
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12307__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _03217_ _03271_ _05563_ _05627_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__and4_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ _02645_ _02693_ _02697_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__a21o_1
XFILLER_5_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5820_ MuI._1462_ MuI._1555_ MuI._1644_ vssd1 vssd1 vccd1 vccd1 MuI._1645_ sky130_fd_sc_hd__o21ai_1
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12247_ _06429_ _04983_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nand2_1
XAuI.pe._700_ AuI.pe._386_ AuI.pe._025_ AuI.pe._078_ AuI.pe.significand\[13\] AuI.pe._036_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._247_ sky130_fd_sc_hd__a221o_1
XMuI._5751_ MuI._1500_ MuI._1502_ MuI._1568_ vssd1 vssd1 vccd1 vccd1 MuI._1569_ sky130_fd_sc_hd__a21o_1
XANTENNA_output70_A net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1625_ AuI._0258_ AuI._0788_ vssd1 vssd1 vccd1 vccd1 AuI._0792_ sky130_fd_sc_hd__or2_1
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12178_ _00555_ _02743_ _02848_ _04011_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a221o_1
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._631_ AuI.pe._029_ AuI.pe._164_ AuI.pe._177_ AuI.pe._182_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._183_ sky130_fd_sc_hd__a211o_1
XFILLER_96_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4702_ MuI._0412_ MuI._0413_ vssd1 vssd1 vccd1 vccd1 MuI._0415_ sky130_fd_sc_hd__nor2_1
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5682_ MuI._2649_ MuI._3246_ MuI._0305_ MuI._2704_ vssd1 vssd1 vccd1 vccd1 MuI._1493_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1556_ AuI._0606_ AuI._0734_ AuI._0735_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[6\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11129_ _03761_ _03769_ _03768_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21o_1
XFILLER_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07781__D _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4633_ MuI._0336_ MuI._0338_ vssd1 vssd1 vccd1 vccd1 MuI._0340_ sky130_fd_sc_hd__nand2_1
XANTENNA__13301__A1 _02705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._562_ AuI.pe.significand\[13\] AuI.pe._383_ AuI.pe._387_ AuI.pe._117_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._118_ sky130_fd_sc_hd__and4_1
XFILLER_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07136__A _06436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1487_ AuI._0629_ AuI._0644_ AuI._0669_ AuI._0672_ vssd1 vssd1 vccd1 vccd1 AuI._0673_
+ sky130_fd_sc_hd__a31o_1
XFILLER_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12977__A _02980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._493_ AuI.pe._033_ vssd1 vssd1 vccd1 vccd1 AuI.pe._055_ sky130_fd_sc_hd__buf_2
XANTENNA_AuI._0907__A1 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4564_ MuI._0209_ MuI._0261_ MuI._0263_ vssd1 vssd1 vccd1 vccd1 MuI._0264_ sky130_fd_sc_hd__a21boi_1
XFILLER_76_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3515_ MuI._1010_ vssd1 vssd1 vccd1 vccd1 MuI._1021_ sky130_fd_sc_hd__buf_4
XMuI._6303_ MuI._2109_ MuI._2113_ vssd1 vssd1 vccd1 vccd1 MuI._2177_ sky130_fd_sc_hd__nor2_1
XANTENNA__09351__A _06544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4495_ MuI._0184_ MuI._0186_ MuI._0187_ vssd1 vssd1 vccd1 vccd1 MuI._0188_ sky130_fd_sc_hd__o21ba_1
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4904__A MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6234_ MuI._2083_ MuI._2100_ vssd1 vssd1 vccd1 vccd1 MuI._2101_ sky130_fd_sc_hd__or2b_1
XANTENNA__06694__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3446_ MuI.a_operand\[25\] MuI.b_operand\[25\] vssd1 vssd1 vccd1 vccd1 MuI._0262_
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09070__B _06611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11615__A1 _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _06460_ _05241_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__nand2_1
XFILLER_205_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11615__B2 _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6165_ MuI._2007_ MuI._2012_ MuI._2017_ vssd1 vssd1 vccd1 vccd1 MuI._2025_ sky130_fd_sc_hd__or3_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08271_ _00882_ _00887_ _00888_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__nand3_1
XFILLER_178_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5116_ MuI._0869_ MuI._0870_ vssd1 vssd1 vccd1 vccd1 MuI._0871_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6096_ MuI._1947_ MuI._1948_ vssd1 vssd1 vccd1 vccd1 MuI._1949_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07222_ _06514_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__nor2_1
XANTENNA__08117__D _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5047_ MuI._0794_ vssd1 vssd1 vccd1 vccd1 MuI._0795_ sky130_fd_sc_hd__inv_2
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07153_ _06447_ _06445_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__and2b_1
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11121__A _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._5706__A1 MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5706__B2 MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _06316_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._0843__B1 net111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08547__A1 _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__A2 _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5949_ MuI._1785_ MuI._1784_ MuI._1783_ MuI._0763_ vssd1 vssd1 vccd1 vccd1 MuI._1787_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11775__B _00197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout114 net52 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout125 net31 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_4
XFILLER_87_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._829_ AuI.operand_a\[28\] AuI.pe._363_ AuI.pe._365_ vssd1 vssd1 vccd1 vccd1
+ AuI.exponent_sub\[5\] sky130_fd_sc_hd__a21bo_1
XFILLER_102_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13048__A _03497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08787__D _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07986_ _00125_ _06433_ _04176_ _00299_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XANTENNA__07691__D _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4142__B1 MuI._2830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07046__A _05917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ _02367_ _02369_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__xor2_1
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06937_ _04747_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[12\] sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_MuI._4086__A MuI.a_operand\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__B1 _00423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4517__C MuI._2790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09656_ _06488_ _04229_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nand2_1
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11854__A1 _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ _04004_ _03690_ _03766_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__and3_1
XANTENNA__06885__A _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__B2 _05895_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08607_ _00991_ _01223_ _01219_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__and3_1
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09587_ _06545_ _04186_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a31o_1
XFILLER_103_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06799_ net51 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__buf_2
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4996__A2 MuI._0421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08538_ _01137_ _01155_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _01084_ _01085_ _01086_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__o21bai_1
XFILLER_23_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _03163_ _04843_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__and2_1
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11480_ _03525_ _04596_ _04099_ _04098_ _04725_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__a32o_1
X_10431_ _02770_ _02928_ _03128_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__or3_1
XFILLER_183_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _06050_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _03054_ _03052_ _03053_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__nand3_1
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ _04926_ _04925_ _04924_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a21bo_1
X_10293_ _00278_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__buf_4
X_13081_ _05900_ _05902_ _05905_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__o21a_1
XANTENNA__08978__C net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _04851_ _04852_ _04816_ _04698_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__o211ai_1
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08340__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1410_ AuI._0139_ vssd1 vssd1 vccd1 vccd1 AuI._0599_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6195__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1341_ AuI._0528_ AuI._0534_ AuI._0535_ vssd1 vssd1 vccd1 vccd1 AuI._0536_ sky130_fd_sc_hd__a21bo_1
XANTENNA_MuI._3612__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12012__D _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ _05785_ _05786_ _05821_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__nor3_1
XAuI._1272_ AuI._0438_ AuI._0350_ vssd1 vssd1 vccd1 vccd1 AuI._0472_ sky130_fd_sc_hd__or2_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07933__A2_N _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06795__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12865_ _05348_ _05482_ _05567_ _05667_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__and4_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4280_ MuI._3340_ MuI._3341_ MuI._3379_ vssd1 vssd1 vccd1 vccd1 MuI._3380_ sky130_fd_sc_hd__and3b_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__A _00077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11816_ _04622_ _02571_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__xnor2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _02741_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and3_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _04545_ _04546_ _04381_ vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__a21oi_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13421__A _05788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _04426_ _04427_ _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a22oi_2
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _06296_ _06299_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__and2b_1
X_10629_ _03341_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__nor2_1
XANTENNA__08234__B _02647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ _02677_ _06209_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_1
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XAuI._0987_ AuI._0163_ vssd1 vssd1 vccd1 vccd1 AuI._0199_ sky130_fd_sc_hd__clkbuf_2
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6852_ MuI._2729_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2758_ sky130_fd_sc_hd__and2b_1
XFILLER_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _06185_ _06186_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__and2_1
XFILLER_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4372__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5803_ MuI._1536_ MuI._1597_ MuI._1624_ MuI._1625_ vssd1 vssd1 vccd1 vccd1 MuI._1627_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3995_ MuI._2517_ MuI._2916_ MuI._2627_ MuI._1318_ vssd1 vssd1 vccd1 vccd1 MuI._3095_
+ sky130_fd_sc_hd__a22o_1
XMuI._6783_ MuI._2685_ MuI._2703_ vssd1 vssd1 vccd1 vccd1 MuI._2705_ sky130_fd_sc_hd__nand2_1
XFILLER_97_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5734_ MuI._1547_ MuI._1548_ MuI._1057_ MuI._1465_ vssd1 vssd1 vccd1 vccd1 MuI._1551_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07201__A1 _06500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1608_ AuI._0708_ AuI._0772_ AuI._0777_ AuI._0778_ vssd1 vssd1 vccd1 vccd1 AuI.result\[15\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07201__B2 _06501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _00036_ _00230_ _00457_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__a21bo_1
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI.pe._614_ AuI.pe._145_ AuI.pe._158_ AuI.pe._141_ vssd1 vssd1 vccd1 vccd1 AuI.pe._167_
+ sky130_fd_sc_hd__or3_1
XFILLER_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._408__D AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5665_ MuI._1473_ MuI._1474_ vssd1 vssd1 vccd1 vccd1 MuI._1475_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._3522__B MuI._0460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._1539_ AuI.pe.Significand\[3\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0722_
+ sky130_fd_sc_hd__or2_1
X_07771_ _00380_ _00381_ _00388_ vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__nand3_1
XFILLER_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._545_ AuI.pe._084_ AuI.pe._070_ AuI.pe._102_ vssd1 vssd1 vccd1 vccd1 AuI.pe._103_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4616_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._0321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09510_ _02120_ _02123_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a211o_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5596_ MuI._1359_ MuI._1358_ MuI._1343_ vssd1 vssd1 vccd1 vccd1 MuI._1399_ sky130_fd_sc_hd__o21ai_1
X_06722_ _02431_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__buf_4
XANTENNA_AuI._1002__A0 net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A1 _04671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__B2 _03306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4547_ MuI._0244_ vssd1 vssd1 vccd1 vccd1 MuI._0245_ sky130_fd_sc_hd__clkbuf_4
XAuI.pe._476_ AuI.pe.significand\[22\] AuI.pe._005_ AuI.pe.significand\[21\] vssd1
+ vssd1 vccd1 vccd1 AuI.pe._040_ sky130_fd_sc_hd__and3b_1
X_09441_ net68 net38 net127 net126 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__and4_1
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4478_ MuI._2671_ MuI._0168_ vssd1 vssd1 vccd1 vccd1 MuI._0169_ sky130_fd_sc_hd__nand2_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4978__A2 MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _01985_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6217_ MuI._2076_ MuI._2080_ MuI._2081_ vssd1 vssd1 vccd1 vccd1 MuI._2082_ sky130_fd_sc_hd__a21bo_1
XMuI._3429_ MuI._0065_ vssd1 vssd1 vccd1 vccd1 MuI.Exception sky130_fd_sc_hd__buf_2
XFILLER_80_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__A1 _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10377__D _00163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ _00933_ _00936_ _00939_ _00940_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__a211o_1
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6148_ MuI.a_operand\[22\] MuI._2693_ MuI._2638_ vssd1 vssd1 vccd1 vccd1 MuI._2006_
+ sky130_fd_sc_hd__and3_1
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10811__A2 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _00641_ _00642_ _00561_ _00643_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6079_ MuI._1894_ MuI._1896_ MuI._1895_ vssd1 vssd1 vccd1 vccd1 MuI._1930_ sky130_fd_sc_hd__o21ba_1
X_07205_ _06502_ _06505_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__nor2_1
XANTENNA__12013__A1 _00270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08185_ _00801_ _00802_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__xnor2_1
XFILLER_119_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07686__D _00303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07136_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__buf_4
XFILLER_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11772__B1 _05112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _06140_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08798__C _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_AuI._1241__A0 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4974__A1_N MuI._1263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ _00335_ _00336_ _00338_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09708_ _02334_ _04100_ _00271_ _01332_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a22o_1
XANTENNA__11827__A1 _02752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ _00345_ _00059_ _03717_ _03718_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nand4_1
XFILLER_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10849__B _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _06560_ _03873_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__nand2_1
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09422__C net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4544__A MuI._2826_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _02965_ _05262_ _05427_ _05426_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a31o_1
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11601_ _00221_ _05520_ _04387_ _04388_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nand4_1
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12581_ _03497_ _05391_ _05314_ _05313_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__a31o_1
XANTENNA__12170__B1_N _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13241__A _03400_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ _04150_ _04152_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__and2_1
XFILLER_211_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._156_ FuI.a_operand\[26\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0910_ net60 net28 vssd1 vssd1 vccd1 vccd1 AuI._0129_ sky130_fd_sc_hd__or2b_1
XFILLER_156_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _04239_ _04237_ _04238_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nand3_1
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFuI._087_ FuI._035_ FuI._043_ FuI._045_ FuI._048_ vssd1 vssd1 vccd1 vccd1 FuI._050_
+ sky130_fd_sc_hd__or4_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _03626_ _05842_ _05906_ _03561_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__a22oi_1
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _02954_ _03112_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__xnor2_4
XANTENNA_MuI._3607__B MuI._0625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._0841_ net111 AuI._0057_ AuI._0058_ AuI._0059_ AuI._0060_ vssd1 vssd1 vccd1 vccd1
+ AuI._0061_ sky130_fd_sc_hd__a221o_1
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _02496_ _04391_ _02743_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__and3_1
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13133_ _03507_ _05842_ _05941_ _05942_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a31o_1
XFILLER_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _03037_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__nor3_1
XFILLER_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09708__B1 _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _05886_ _05955_ _05960_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__or3_1
XANTENNA__10318__A1 _02959_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ _02962_ _02963_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__nor2_1
XANTENNA__10318__B2 _00217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XMuI._3780_ MuI.b_operand\[3\] vssd1 vssd1 vccd1 vccd1 MuI._2880_ sky130_fd_sc_hd__buf_2
X_12015_ _03378_ _00279_ _05187_ _05252_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nand4_2
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0854__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5450_ MuI._1178_ MuI._1237_ vssd1 vssd1 vccd1 vccd1 MuI._1238_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1324_ AuI._0257_ AuI._0517_ AuI._0518_ AuI._0519_ vssd1 vssd1 vccd1 vccd1 AuI._0521_
+ sky130_fd_sc_hd__a31oi_2
XFILLER_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4401_ MuI._0081_ MuI._0083_ vssd1 vssd1 vccd1 vccd1 MuI._0084_ sky130_fd_sc_hd__or2b_1
XANTENNA__09487__A2 _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5381_ MuI._1158_ MuI._1159_ MuI._1160_ vssd1 vssd1 vccd1 vccd1 MuI._1162_ sky130_fd_sc_hd__and3_1
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07414__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07498__A1 _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ _03550_ _03615_ _05585_ _05649_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__and4_1
XAuI._1255_ AuI._0455_ AuI._0456_ vssd1 vssd1 vccd1 vccd1 AuI._0457_ sky130_fd_sc_hd__and2_1
XFILLER_62_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3880__A2 MuI._2850_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4332_ MuI._0006_ MuI._0008_ vssd1 vssd1 vccd1 vccd1 MuI._0009_ sky130_fd_sc_hd__xor2_1
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _05712_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__xnor2_1
XAuI._1186_ AuI._0261_ AuI._0388_ AuI._0391_ vssd1 vssd1 vccd1 vccd1 AuI._0392_ sky130_fd_sc_hd__nand3_4
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI.pe._475__A1 AuI.pe._013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4263_ MuI._3362_ vssd1 vssd1 vccd1 vccd1 MuI._3363_ sky130_fd_sc_hd__clkbuf_4
XMuI._6002_ MuI._3111_ MuI._3117_ MuI._1844_ vssd1 vssd1 vccd1 vccd1 MuI._1845_ sky130_fd_sc_hd__a21oi_2
X_12779_ _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__or2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4194_ MuI._3292_ MuI._3293_ vssd1 vssd1 vccd1 vccd1 MuI._3294_ sky130_fd_sc_hd__and2_1
XANTENNA__10254__B1 _02741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10494__B _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _01311_ _01312_ _01313_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__o21ai_1
XFILLER_131_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6835_ MuI._2724_ MuI._2737_ vssd1 vssd1 vccd1 vccd1 MuI._2750_ sky130_fd_sc_hd__and2b_1
XFILLER_103_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _01556_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6766_ MuI._2608_ MuI._2612_ vssd1 vssd1 vccd1 vccd1 MuI._2686_ sky130_fd_sc_hd__or2_1
XFILLER_97_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3978_ MuI._3075_ MuI._3076_ vssd1 vssd1 vccd1 vccd1 MuI._3078_ sky130_fd_sc_hd__xnor2_1
X_08872_ _01488_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__nor2_1
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5717_ MuI._1525_ MuI._1530_ MuI._1531_ vssd1 vssd1 vccd1 vccd1 MuI._1532_ sky130_fd_sc_hd__nand3_1
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07823_ _00440_ _00247_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__nor2_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6697_ MuI._2602_ MuI._2609_ vssd1 vssd1 vccd1 vccd1 MuI._2610_ sky130_fd_sc_hd__or2_1
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5648_ MuI._1242_ MuI._1455_ vssd1 vssd1 vccd1 vccd1 MuI._1456_ sky130_fd_sc_hd__xor2_1
X_07754_ _00186_ _00187_ _00209_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__nor3_1
XAuI.pe._528_ AuI.pe._014_ AuI.pe._086_ AuI.pe._066_ AuI.pe._033_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._087_ sky130_fd_sc_hd__a22o_1
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06705_ _02248_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__clkbuf_8
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5579_ MuI._2882_ MuI._0320_ vssd1 vssd1 vccd1 vccd1 MuI._1380_ sky130_fd_sc_hd__nand2_1
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07685_ _06433_ vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._459_ AuI.pe.significand\[24\] vssd1 vssd1 vccd1 vccd1 AuI.pe._024_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08139__B _06579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09424_ _02043_ _02044_ _06544_ _00074_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10493__B1 _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5179__B MuI._0320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09355_ net111 _04574_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__nand2_1
XANTENNA__13431__B1 _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13061__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _00920_ _00922_ _00923_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__o21bai_1
X_09286_ _01787_ _01786_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__and2b_1
XANTENNA__08155__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _00852_ _00853_ _00854_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__or3_1
XANTENNA__07994__A _00610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__C1 _05992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08305__D _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08168_ _06501_ _06500_ _05756_ _00785_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__and4_1
XANTENNA__07950__A1_N _03002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ _06423_ vssd1 vssd1 vccd1 vccd1 FuI.a_operand\[28\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08099_ _00221_ _04918_ _00715_ _00716_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__nand4_1
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__B _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ _03239_ _05338_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__and2b_1
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _03928_ _02728_ _02732_ AuI.result\[0\] vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09714__A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09433__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09469__A2 _00035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10579__B _03289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07234__A _06534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ _03700_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__xor2_4
XANTENNA__08049__B _00519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _02614_ _02609_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or2_1
XAuI._1040_ AuI._0251_ vssd1 vssd1 vccd1 vccd1 AuI._0252_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _03625_ _03627_ _03445_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a21o_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12633_ _05495_ _05497_ _05493_ _05494_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__a211o_1
XFILLER_169_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ _06434_ _00678_ _00412_ _00530_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and4_1
XFILLER_200_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5367__A2 MuI._0305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _04094_ _04183_ _04296_ _04297_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a211oi_4
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12495_ _04997_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__inv_2
XFuI._139_ FuI._001_ net145 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[10\] sky130_fd_sc_hd__dlxtn_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11446_ _04220_ _04221_ _04067_ _04187_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__o211ai_2
XFILLER_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4866__A1_N MuI._2841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4950_ MuI._0682_ MuI._0687_ vssd1 vssd1 vccd1 vccd1 MuI._0688_ sky130_fd_sc_hd__and2_1
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XAuI._0824_ net44 vssd1 vssd1 vccd1 vccd1 AuI._0044_ sky130_fd_sc_hd__inv_2
XFILLER_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _04025_ _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3901_ MuI._2754_ MuI._2605_ MuI._2660_ MuI._3000_ vssd1 vssd1 vccd1 vccd1 MuI._3001_
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07955__A2 _00085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13116_ _03561_ _05842_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__nand2_1
XANTENNA_MuI._5552__B MuI._0445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4881_ MuI._0524_ MuI._0525_ MuI._0527_ MuI._0491_ vssd1 vssd1 vccd1 vccd1 MuI._0612_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10328_ _03016_ _03017_ _03018_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__a21oi_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6620_ MuI._2523_ MuI._2524_ vssd1 vssd1 vccd1 vccd1 MuI._2525_ sky130_fd_sc_hd__nor2_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._3832_ MuI._2682_ MuI._2930_ MuI._2931_ vssd1 vssd1 vccd1 vccd1 MuI._2932_ sky130_fd_sc_hd__a21bo_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__inv_2
X_10259_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12161__B1 _04991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3763_ MuI._2861_ MuI._2862_ vssd1 vssd1 vccd1 vccd1 MuI._2863_ sky130_fd_sc_hd__xnor2_1
XMuI._6551_ MuI._2232_ MuI._2448_ vssd1 vssd1 vccd1 vccd1 MuI._2449_ sky130_fd_sc_hd__and2_1
XFILLER_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5502_ MuI._1258_ MuI._1249_ MuI._1257_ vssd1 vssd1 vccd1 vccd1 MuI._1295_ sky130_fd_sc_hd__nand3_1
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6482_ MuI._1922_ MuI._1921_ vssd1 vssd1 vccd1 vccd1 MuI._2373_ sky130_fd_sc_hd__or2b_1
XMuI._3694_ MuI._1274_ MuI._2787_ MuI._2793_ MuI._2788_ vssd1 vssd1 vccd1 vccd1 MuI._2794_
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5433_ MuI._1211_ MuI._1206_ vssd1 vssd1 vccd1 vccd1 MuI._1220_ sky130_fd_sc_hd__or2b_1
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1307_ AuI._0503_ AuI._0504_ AuI._0486_ vssd1 vssd1 vccd1 vccd1 AuI._0505_ sky130_fd_sc_hd__or3b_1
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3800__B MuI._0768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5364_ MuI._1141_ MuI._1143_ vssd1 vssd1 vccd1 vccd1 MuI._1144_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07470_ net49 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__buf_6
XAuI._1238_ AuI._0420_ AuI._0425_ AuI._0440_ vssd1 vssd1 vccd1 vccd1 AuI._0441_ sky130_fd_sc_hd__a21o_1
XANTENNA__06983__A _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4315_ MuI._3261_ MuI._3414_ vssd1 vssd1 vccd1 vccd1 MuI._3415_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5295_ MuI._2885_ MuI._3362_ MuI._2881_ MuI._0085_ vssd1 vssd1 vccd1 vccd1 MuI._1068_
+ sky130_fd_sc_hd__a22o_1
XAuI._1169_ AuI._0370_ AuI._0372_ AuI._0375_ AuI._0288_ AuI._0249_ vssd1 vssd1 vccd1
+ vccd1 AuI._0376_ sky130_fd_sc_hd__a221oi_4
XFILLER_195_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4246_ MuI._2473_ MuI._2363_ vssd1 vssd1 vccd1 vccd1 MuI._3346_ sky130_fd_sc_hd__nand2_1
X_09140_ _01736_ _01755_ _01756_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or4b_2
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11975__B1 _05638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12209__B _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4177_ MuI._3165_ MuI._3275_ MuI._3258_ vssd1 vssd1 vccd1 vccd1 MuI._3277_ sky130_fd_sc_hd__and3_1
XFILLER_175_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3528__A MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ _06491_ _06602_ _06604_ _06492_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08840__B1 _06581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08022_ _06511_ _06512_ _06532_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__and3_1
XFILLER_175_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4030__A2 MuI._2975_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__A1_N _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07319__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09973_ _02634_ _02637_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__nand2_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6818_ MuI._2712_ MuI._2738_ vssd1 vssd1 vccd1 vccd1 MuI._2740_ sky130_fd_sc_hd__and2b_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08924_ _01541_ _01217_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__xnor2_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4078__B MuI._3158_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6749_ MuI._1747_ MuI._2308_ MuI._2475_ MuI._2477_ vssd1 vssd1 vccd1 vccd1 MuI._2667_
+ sky130_fd_sc_hd__o31a_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08855_ _01462_ _01463_ _01464_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__o21ba_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ _02808_ _00423_ _00002_ _02765_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a22oi_2
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09253__B _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _01402_ _01388_ _01393_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__and3_1
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _00350_ _00352_ _00351_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__a21o_1
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06893__A _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _00268_ _00273_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._6243__B1 MuI._1483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07204__D _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__B1 _06591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _02024_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nor2_1
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4244__D MuI._2495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07599_ _00028_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__buf_4
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11304__A _03228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09338_ _01840_ _01925_ _01955_ _01952_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__o211a_1
XFILLER_139_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09269_ _06479_ _06480_ net6 net7 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__and4_1
XFILLER_138_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ _03955_ _03954_ _03953_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__a21bo_1
XFILLER_193_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12280_ _05118_ _05119_ _05037_ _04984_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__a211oi_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _03904_ _03905_ _03989_ _03990_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a22o_1
XFILLER_181_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11162_ _03912_ _03915_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nor2_1
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__inv_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11093_ _02388_ _04262_ _02743_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__and3_1
XFILLER_95_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13486__A3 _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A a_operand[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _03906_ _02118_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__nand2b_2
XANTENNA__07890__C _06431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11249__A2 _01988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10102__B _05402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ _04740_ _04742_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__nand2_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10946_ _02883_ _03322_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__and2b_1
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1023_ AuI._0209_ AuI._0222_ AuI._0234_ AuI._0152_ vssd1 vssd1 vccd1 vccd1 AuI._0235_
+ sky130_fd_sc_hd__a211o_1
XFILLER_205_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4100_ MuI._2840_ MuI._2605_ MuI._2836_ MuI._2854_ vssd1 vssd1 vccd1 vccd1 MuI._3200_
+ sky130_fd_sc_hd__and4_1
X_10877_ _03606_ _03607_ _03608_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5080_ MuI._0829_ MuI._0830_ MuI._2850_ MuI.a_operand\[0\] vssd1 vssd1 vccd1
+ vccd1 MuI._0831_ sky130_fd_sc_hd__and4bb_1
XANTENNA__11214__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _05348_ _05359_ _05346_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a21o_1
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4031_ MuI._3128_ MuI._3129_ MuI._3130_ vssd1 vssd1 vccd1 vccd1 MuI._3131_ sky130_fd_sc_hd__nand3b_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ _03174_ _03257_ _05406_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__nand4_1
XANTENNA__08822__B1 _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11868__B _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4012__A2 MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _05289_ _05290_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a22oi_2
XANTENNA__08523__A _00915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5982_ MuI._1819_ MuI._1821_ vssd1 vssd1 vccd1 vccd1 MuI._1823_ sky130_fd_sc_hd__and2_1
X_11429_ _03324_ _05047_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nand2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__C _00385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6378__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4933_ MuI._0667_ MuI._0668_ vssd1 vssd1 vccd1 vccd1 MuI._0670_ sky130_fd_sc_hd__nand2_1
XFILLER_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0807_ net17 vssd1 vssd1 vccd1 vccd1 AuI._0027_ sky130_fd_sc_hd__inv_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._5713__D MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._793_ AuI.pe._332_ vssd1 vssd1 vccd1 vccd1 AuI.pe._333_ sky130_fd_sc_hd__inv_2
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4864_ MuI._0591_ MuI._0593_ MuI._2841_ MuI._2352_ vssd1 vssd1 vccd1 vccd1 MuI._0594_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06970_ _05101_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__buf_4
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06978__A _05187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6603_ MuI._1836_ MuI._1839_ vssd1 vssd1 vccd1 vccd1 MuI._2507_ sky130_fd_sc_hd__and2b_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3815_ MuI._2860_ MuI._2914_ vssd1 vssd1 vccd1 vccd1 MuI._2915_ sky130_fd_sc_hd__nand2_1
XANTENNA__08896__C _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4795_ MuI._0510_ MuI._0514_ MuI._0516_ vssd1 vssd1 vccd1 vccd1 MuI._0518_ sky130_fd_sc_hd__or3_1
XFILLER_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06697__B _02053_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6534_ MuI._2221_ MuI._2222_ MuI._2219_ vssd1 vssd1 vccd1 vccd1 MuI._2431_ sky130_fd_sc_hd__o21bai_1
XMuI._3746_ MuI._2843_ MuI._2844_ MuI._2845_ MuI._1472_ vssd1 vssd1 vccd1 vccd1 MuI._2846_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08640_ _01256_ _01257_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__nand2_1
XFILLER_26_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6465_ MuI._2315_ MuI._2316_ MuI._2317_ vssd1 vssd1 vccd1 vccd1 MuI._2355_ sky130_fd_sc_hd__o21ai_1
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3677_ MuI._2765_ vssd1 vssd1 vccd1 vccd1 MuI._2773_ sky130_fd_sc_hd__clkbuf_4
X_08571_ _01156_ _01172_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__or2_1
XFILLER_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5416_ MuI._1191_ MuI._1199_ MuI._1200_ vssd1 vssd1 vccd1 vccd1 MuI._1201_ sky130_fd_sc_hd__a21bo_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _00138_ _00139_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__and2b_1
XMuI._6396_ MuI._2274_ MuI._2277_ MuI._2251_ MuI._2267_ vssd1 vssd1 vccd1 vccd1 MuI._2279_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5347_ MuI._3363_ MuI._3185_ MuI._0101_ MuI._2892_ vssd1 vssd1 vccd1 vccd1 MuI._1125_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__07602__A _03013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07453_ _00044_ _00055_ _00068_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__and3_1
XANTENNA__13323__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10666__C _00002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._5278_ MuI._1046_ MuI._1047_ MuI._1030_ vssd1 vssd1 vccd1 vccd1 MuI._1049_ sky130_fd_sc_hd__a21o_1
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5457__B MuI._3307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ _06517_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__buf_4
XFILLER_50_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4251__A2 MuI._2786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._1295__D AuI._0493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._4229_ MuI._3326_ MuI._3327_ MuI._3328_ vssd1 vssd1 vccd1 vccd1 MuI._3329_ sky130_fd_sc_hd__o21ba_1
XFILLER_124_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _00221_ _03873_ _01424_ _01425_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _01665_ _01666_ _01671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__nor3b_2
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07975__C _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09369__A1 _02474_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ _06496_ _06490_ _06493_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__or3_1
XANTENNA__09369__B2 _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07049__A _05948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _02608_ _02613_ _02619_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__and3b_1
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06888__A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08907_ _06610_ _04316_ _01522_ _01523_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__o2bb2a_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _02516_ _02526_ _02530_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or4bb_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08838_ _01444_ _01443_ _01442_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._4536__B MuI._3372_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _01383_ _01386_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__xnor2_2
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10800_ _03524_ _03526_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__xor2_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _04581_ _04579_ _04580_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__nand3_2
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07512__A _00086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A2_N _04186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _03450_ _03451_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nand3b_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _06170_ _06342_ _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ _03195_ _03214_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__nand2_1
XFILLER_201_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ MuI.result\[15\] _02738_ _04642_ _04865_ _05250_ vssd1 vssd1 vccd1 vccd1
+ _05251_ sky130_fd_sc_hd__a221o_1
XANTENNA__10295__D _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _06292_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__or2_1
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10593_ _02720_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ _05174_ _05175_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__or2_1
XFILLER_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09158__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _05099_ _05100_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a21o_1
XFILLER_123_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _00086_ _06623_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__and2_2
XAuI._1641_ AuI._0804_ vssd1 vssd1 vccd1 vccd1 AuI.result\[22\] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ _02848_ _05003_ _00555_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__a21o_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 ALU_Output[13] sky130_fd_sc_hd__buf_2
XFILLER_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11145_ _03896_ _03897_ _03727_ _03880_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a211o_1
XANTENNA__12015__D _05252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 ALU_Output[23] sky130_fd_sc_hd__buf_2
XAuI._1572_ AuI._0606_ AuI._0747_ AuI._0748_ AuI._0700_ vssd1 vssd1 vccd1 vccd1 AuI.result\[9\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 ALU_Output[4] sky130_fd_sc_hd__buf_2
XFILLER_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11076_ _03647_ _03649_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__nand2_1
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3600_ MuI._0889_ MuI._1043_ MuI._1945_ vssd1 vssd1 vccd1 vccd1 MuI._1956_ sky130_fd_sc_hd__and3_1
XMuI._4580_ MuI._0275_ MuI._0276_ MuI._0280_ vssd1 vssd1 vccd1 vccd1 MuI._0281_ sky130_fd_sc_hd__a21boi_1
X_10027_ _02685_ _02687_ _02690_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__o21a_1
XANTENNA__11209__A _00133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3531_ MuI._1175_ MuI._1186_ vssd1 vssd1 vccd1 vccd1 MuI._1197_ sky130_fd_sc_hd__nor2_1
XANTENNA__12419__A1 _01146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__B2 _01147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0862__A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6250_ MuI._2115_ MuI._2116_ vssd1 vssd1 vccd1 vccd1 MuI._2118_ sky130_fd_sc_hd__nor2_1
XMuI._3462_ MuI._0427_ vssd1 vssd1 vccd1 vccd1 MuI._0438_ sky130_fd_sc_hd__clkbuf_2
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11978_ _04793_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__or3_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5201_ MuI._0960_ MuI._0954_ MuI._0956_ vssd1 vssd1 vccd1 vccd1 MuI._0964_ sky130_fd_sc_hd__nand3_1
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._6181_ MuI._2034_ MuI._2041_ vssd1 vssd1 vccd1 vccd1 MuI._2042_ sky130_fd_sc_hd__nand2_1
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07422__A _04703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ _03660_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__nand2_1
XFILLER_189_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5132_ MuI._2873_ MuI._3190_ MuI._0085_ MuI.a_operand\[6\] vssd1 vssd1 vccd1
+ vccd1 MuI._0888_ sky130_fd_sc_hd__and4_1
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI._1006_ net120 net11 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0218_ sky130_fd_sc_hd__mux2_1
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MuI._4181__B MuI._3279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5063_ MuI._0799_ MuI._0805_ vssd1 vssd1 vccd1 vccd1 MuI._0813_ sky130_fd_sc_hd__xnor2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4014_ MuI._0361_ MuI._0603_ MuI._2791_ MuI._2787_ vssd1 vssd1 vccd1 vccd1 MuI._3114_
+ sky130_fd_sc_hd__and4_1
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3992__A1 MuI._3091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09349__A _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5965_ MuI._1801_ MuI._1803_ MuI._1798_ vssd1 vssd1 vccd1 vccd1 MuI._1805_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4916_ MuI._0633_ MuI._0646_ MuI._0649_ MuI._0650_ vssd1 vssd1 vccd1 vccd1 MuI._0651_
+ sky130_fd_sc_hd__o211ai_2
XFILLER_114_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ _06469_ _00150_ net126 net125 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__and4_1
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5896_ MuI._0727_ MuI._1724_ MuI._1726_ MuI._1728_ vssd1 vssd1 vccd1 vccd1 MuI._1729_
+ sky130_fd_sc_hd__nor4_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4847_ MuI._0327_ MuI._3189_ MuI._3190_ MuI._2429_ vssd1 vssd1 vccd1 vccd1 MuI._0575_
+ sky130_fd_sc_hd__a22oi_1
X_09741_ _02376_ _02384_ _02385_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__o211ai_4
XANTENNA__09084__A _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06953_ _04918_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12222__B _00132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4778_ MuI._0312_ MuI._0498_ vssd1 vssd1 vccd1 vccd1 MuI._0499_ sky130_fd_sc_hd__nor2_1
X_09672_ _02263_ _02288_ _02309_ _02312_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a211o_1
XFILLER_95_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06884_ _04176_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__buf_4
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6517_ MuI._2132_ MuI._1780_ vssd1 vssd1 vccd1 vccd1 MuI._2412_ sky130_fd_sc_hd__and2b_1
XMuI._3729_ MuI.a_operand\[5\] vssd1 vssd1 vccd1 vccd1 MuI._2829_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08623_ _01034_ _01227_ _01226_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__a21o_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10958__A _03534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6448_ MuI._2333_ MuI._2335_ vssd1 vssd1 vccd1 vccd1 MuI._2336_ sky130_fd_sc_hd__and2_1
XANTENNA_AuI.pe._443__B AuI.pe.significand\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _01157_ _01171_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__nand2_1
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07332__A _06598_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _00077_ _04316_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__nand2_2
XFILLER_211_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6379_ MuI._2258_ MuI._2259_ vssd1 vssd1 vccd1 vccd1 MuI._2260_ sky130_fd_sc_hd__nor2_1
XANTENNA__11094__B1 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08485_ _01098_ _01102_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07436_ _00042_ _00053_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4091__B MuI._1461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07367_ _06664_ _06665_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__nand3b_1
XFILLER_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _01697_ _01700_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__nand2_1
XFILLER_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07298_ net41 vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__clkbuf_4
XFILLER_136_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _01210_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__xnor2_2
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0861__B2 net106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11020__C _03762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12897__A1 _03346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__B2 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09762__A1 _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__B2 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__A2_N _00272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__B _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__B_N _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07507__A net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09939_ _02328_ _02588_ _02589_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__and3_1
XANTENNA_MuI._4547__A MuI._0244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12132__B _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__B _06515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _05838_ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nand2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11901_ _04711_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__xor2_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11971__B _03047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _05338_ _02718_ _02721_ _03174_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__a221o_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._4999__B1 MuI._3396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _02871_ _04636_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__or2_1
XANTENNA__09441__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5660__A1 MuI._1813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MuI._5660__B2 MuI._1318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__A1 _00046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _04563_ _04564_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__xor2_4
XFILLER_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07828__B2 _00049_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _03423_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__nand3_1
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _02713_ _04346_ _04491_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__o21ai_4
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ _05853_ _02726_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__nor2_1
XANTENNA__11699__A _02860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ _00345_ _04531_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a22o_1
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09169__A _02582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ _06185_ _06244_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__nor2_1
XANTENNA__08907__A2_N _04316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10576_ _03108_ _03111_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nor2_1
XFILLER_182_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12307__B _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ _00231_ _03424_ _00382_ _00299_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a22oi_1
XFILLER_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295_ _02833_ _06146_ _06151_ _06205_ _03489_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o311a_1
XANTENNA_AuI._0852__B2 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__xor2_4
XFILLER_142_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5750_ MuI._1565_ MuI._1567_ vssd1 vssd1 vccd1 vccd1 MuI._1568_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1624_ AuI._0678_ AuI._0684_ vssd1 vssd1 vccd1 vccd1 AuI._0791_ sky130_fd_sc_hd__xor2_1
X_12177_ MuI.result\[13\] _02736_ _02944_ _04736_ vssd1 vssd1 vccd1 vccd1 _05011_
+ sky130_fd_sc_hd__a22o_1
XAuI.pe._630_ AuI.pe._106_ AuI.pe._066_ AuI.pe._178_ AuI.pe._181_ vssd1 vssd1 vccd1
+ vccd1 AuI.pe._182_ sky130_fd_sc_hd__a211o_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12323__A _03163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4701_ MuI._0412_ MuI._0413_ vssd1 vssd1 vccd1 vccd1 MuI._0414_ sky130_fd_sc_hd__xor2_1
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5681_ MuI._2799_ MuI._2918_ MuI._0228_ MuI._3371_ vssd1 vssd1 vccd1 vccd1 MuI._1492_
+ sky130_fd_sc_hd__and4_1
XANTENNA__07417__A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _03543_ _03547_ _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a211oi_1
XAuI._1555_ AuI.pe.Significand\[6\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0735_
+ sky130_fd_sc_hd__or2_1
XFILLER_122_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._561_ AuI.pe.significand\[14\] AuI.pe.significand\[15\] AuI.pe._367_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._117_ sky130_fd_sc_hd__nor3_1
XMuI._4632_ MuI._0210_ MuI._0337_ vssd1 vssd1 vccd1 vccd1 MuI._0338_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11059_ _03623_ _03625_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__nand2_1
XFILLER_37_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1486_ AuI._0670_ AuI._0671_ vssd1 vssd1 vccd1 vccd1 AuI._0672_ sky130_fd_sc_hd__or2_1
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07516__B1 _00048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._492_ AuI.pe._053_ vssd1 vssd1 vccd1 vccd1 AuI.pe._054_ sky130_fd_sc_hd__buf_2
XANTENNA_AuI.pe._544__A AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__B _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4563_ MuI._0206_ MuI._0208_ vssd1 vssd1 vccd1 vccd1 MuI._0263_ sky130_fd_sc_hd__nand2_1
XANTENNA__09632__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6302_ MuI._2173_ MuI._2174_ vssd1 vssd1 vccd1 vccd1 MuI._2175_ sky130_fd_sc_hd__nor2_1
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3514_ MuI.a_operand\[19\] vssd1 vssd1 vccd1 vccd1 MuI._1010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4494_ MuI._2440_ MuI._2844_ MuI._2451_ MuI._2845_ vssd1 vssd1 vccd1 vccd1 MuI._0187_
+ sky130_fd_sc_hd__and4_1
XANTENNA__09351__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6233_ MuI._2083_ MuI._2084_ MuI._2098_ vssd1 vssd1 vccd1 vccd1 MuI._2100_ sky130_fd_sc_hd__or3_1
XANTENNA_MuI._4904__B MuI._0245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3445_ MuI.a_operand\[26\] MuI.b_operand\[26\] vssd1 vssd1 vccd1 vccd1 MuI._0251_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07152__A _03669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__A2 _00530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12993__A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._6164_ MuI._2019_ MuI._2023_ vssd1 vssd1 vccd1 vccd1 MuI._2024_ sky130_fd_sc_hd__or2b_1
XANTENNA_MuI._4623__C MuI._2837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _00574_ _00881_ _00880_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__a21o_1
XANTENNA__06991__A _05327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5115_ MuI._2352_ MuI._2966_ vssd1 vssd1 vccd1 vccd1 MuI._0870_ sky130_fd_sc_hd__nand2_1
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _06514_ _06521_ _02528_ _05112_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and4bb_1
XMuI._6095_ MuI._1864_ MuI._1866_ MuI._1865_ vssd1 vssd1 vccd1 vccd1 MuI._1948_ sky130_fd_sc_hd__o21ba_1
XFILLER_193_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5046_ MuI._2799_ MuI._2918_ MuI.a_operand\[1\] MuI.a_operand\[0\] vssd1 vssd1
+ vccd1 vccd1 MuI._0794_ sky130_fd_sc_hd__and4_1
XFILLER_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07152_ _03669_ _03895_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nand2_1
XFILLER_146_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11121__B _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5706__A2 MuI._2892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _04671_ _06284_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__and2_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._0843__A1 net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12879__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5948_ MuI._0763_ MuI._1783_ MuI._1784_ MuI._1785_ vssd1 vssd1 vccd1 vccd1 MuI._1786_
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__08547__A2 _03884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13329__A _03820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 FuI.a_operand\[24\] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_2
XFILLER_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout115 net5 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._828_ AuI.pe._360_ AuI.pe._362_ AuI.pe._364_ vssd1 vssd1 vccd1 vccd1 AuI.pe._365_
+ sky130_fd_sc_hd__a21o_1
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout126 net30 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5879_ MuI._1649_ MuI._1709_ vssd1 vssd1 vccd1 vccd1 MuI._1710_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13048__B _05831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ _00309_ _00311_ _00310_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__o21ai_1
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XAuI.pe._759_ AuI.pe.significand\[3\] AuI.pe._012_ AuI.pe._300_ AuI.pe._014_ AuI.pe._302_
+ vssd1 vssd1 vccd1 vccd1 AuI.pe._303_ sky130_fd_sc_hd__a221o_1
X_09724_ _02278_ _02368_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06936_ _04736_ _04402_ _04478_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and3_1
XANTENNA__07688__A1_N _00283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11303__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4086__B MuI._2894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11303__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4517__D MuI._3223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _02248_ _04305_ _02247_ _02246_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06867_ _03993_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__buf_4
XANTENNA__11854__A2 _05777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08606_ _00991_ _01219_ _01223_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a21o_1
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09586_ _01332_ _06480_ _00266_ _00592_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__and4_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06798_ _03250_ vssd1 vssd1 vccd1 vccd1 MuI.b_operand\[21\] sky130_fd_sc_hd__clkbuf_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07062__A _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _01153_ _01154_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__nand2_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._4533__C MuI._2829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07997__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _06598_ _06599_ _04509_ _00035_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__and4_1
XFILLER_184_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ _00031_ _00034_ net119 _00036_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__and4bb_1
XFILLER_184_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08399_ _00986_ _01003_ _01015_ _01016_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a211oi_4
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _02770_ _02928_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__o21ai_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MuI._3446__A MuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _03052_ _03053_ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__a21o_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ _04924_ _04925_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__nand3b_1
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _05976_ _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__xnor2_1
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10292_ _02980_ _00093_ _04520_ _00281_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09735__A1 _02604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _04816_ _04698_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a211o_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08978__D net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08340__B _05241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__B1 _00363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6195__C MuI._2849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._1340_ AuI._0526_ AuI._0527_ vssd1 vssd1 vccd1 vccd1 AuI._0535_ sky130_fd_sc_hd__nand2_1
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _05785_ _05786_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__o21a_1
XAuI._1271_ AuI._0330_ AuI._0356_ vssd1 vssd1 vccd1 vccd1 AuI._0471_ sky130_fd_sc_hd__nor2_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12864_ _05746_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and2_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _02572_ _02551_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__or2b_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__B _00550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output101_A net101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ _02596_ _02628_ _05576_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__nand3_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10110__B _02550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _04381_ _04545_ _04546_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__and3_1
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11677_ _04426_ _04427_ _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__and4_1
XANTENNA_AuI._1674__C AuI._0138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13416_ _06328_ _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__or2b_1
X_10628_ _06444_ _00676_ _00090_ _00093_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__and4_1
XFILLER_167_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09423__B1 _04434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._5149__B1 MuI._2881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08234__C _06602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ _02831_ _02830_ _06205_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__or3b_1
XFILLER_127_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ _03091_ _03093_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nor2_1
XAuI._0986_ AuI._0197_ vssd1 vssd1 vccd1 vccd1 AuI._0198_ sky130_fd_sc_hd__inv_2
XANTENNA_AuI._0825__B2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6851_ MuI._2728_ MuI._2757_ vssd1 vssd1 vccd1 vccd1 MuI.result\[19\] sky130_fd_sc_hd__nor2_1
XFILLER_115_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11876__B _04685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13278_ _06185_ _06186_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and3_1
XANTENNA__08531__A _03335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5802_ MuI._1622_ MuI._1623_ MuI._1607_ vssd1 vssd1 vccd1 vccd1 MuI._1625_ sky130_fd_sc_hd__a21oi_1
XANTENNA_MuI._4372__A1 MuI._2440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MuI._4372__B2 MuI._2671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6782_ MuI._2577_ MuI._2580_ MuI._2587_ vssd1 vssd1 vccd1 vccd1 MuI._2703_ sky130_fd_sc_hd__a21o_1
X_12229_ _05056_ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__xnor2_1
XMuI._3994_ MuI._1318_ MuI._1813_ MuI._2916_ MuI._2627_ vssd1 vssd1 vccd1 vccd1 MuI._3094_
+ sky130_fd_sc_hd__nand4_1
XFILLER_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6386__B MuI._2851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5733_ MuI._1057_ MuI._1465_ MuI._1547_ MuI._1548_ vssd1 vssd1 vccd1 vccd1 MuI._1550_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12730__B1 _05884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1607_ AuI.pe.Significand\[15\] AuI._0695_ AuI.Exception vssd1 vssd1 vccd1 vccd1
+ AuI._0778_ sky130_fd_sc_hd__o21ba_1
XFILLER_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07201__A2 _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._613_ AuI.pe._030_ AuI.pe._164_ AuI.pe._112_ AuI.pe._059_ AuI.pe._165_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._166_ sky130_fd_sc_hd__a221o_1
XFILLER_110_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5664_ MuI._0986_ MuI._1471_ vssd1 vssd1 vccd1 vccd1 MuI._1474_ sky130_fd_sc_hd__or2_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1538_ AuI._0599_ vssd1 vssd1 vccd1 vccd1 AuI._0721_ sky130_fd_sc_hd__clkbuf_2
X_07770_ _00383_ _00387_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06986__A _05273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI.pe._544_ AuI.pe._393_ vssd1 vssd1 vccd1 vccd1 AuI.pe._102_ sky130_fd_sc_hd__buf_2
XMuI._4615_ MuI.a_operand\[0\] vssd1 vssd1 vccd1 vccd1 MuI._0320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06721_ _02420_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__buf_4
XMuI._5595_ MuI._1359_ MuI._1343_ MuI._1358_ vssd1 vssd1 vccd1 vccd1 MuI._1398_ sky130_fd_sc_hd__or3_1
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_AuI._1002__A1 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A2 _02941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1469_ AuI._0342_ AuI._0346_ vssd1 vssd1 vccd1 vccd1 AuI._0655_ sky130_fd_sc_hd__and2b_1
XAuI.pe._475_ AuI.pe._013_ AuI.pe._014_ AuI.pe._033_ vssd1 vssd1 vccd1 vccd1 AuI.pe._039_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_65_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4546_ MuI.a_operand\[1\] vssd1 vssd1 vccd1 vccd1 MuI._0244_ sky130_fd_sc_hd__clkbuf_4
X_09440_ _01999_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__nor2_1
XANTENNA__13038__A1 _03293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4477_ MuI.b_operand\[8\] vssd1 vssd1 vccd1 vccd1 MuI._0168_ sky130_fd_sc_hd__buf_2
X_09371_ _01986_ _01987_ _01891_ _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07425__A2_N _00036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__C _01026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6216_ MuI._2038_ MuI._2079_ MuI._2078_ vssd1 vssd1 vccd1 vccd1 MuI._2081_ sky130_fd_sc_hd__nand3_1
XMuI._3428_ MuI.b_operand\[24\] MuI.b_operand\[25\] MuI._0021_ MuI._0054_ vssd1 vssd1
+ vccd1 vccd1 MuI._0065_ sky130_fd_sc_hd__a31o_1
XANTENNA__12797__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _00618_ _00938_ _00937_ _00900_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a211oi_1
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__A2 _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A1 _01071_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6147_ MuI._1996_ MuI._2004_ vssd1 vssd1 vccd1 vccd1 MuI._2005_ sky130_fd_sc_hd__nand2_1
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _00849_ _00868_ _00869_ _00870_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__and4b_2
XFILLER_166_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11132__A _02983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ _06503_ _06504_ _05370_ _05434_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__and4_1
XMuI._6078_ MuI._1285_ MuI._2849_ MuI._1856_ MuI._1854_ vssd1 vssd1 vccd1 vccd1 MuI._1929_
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _00409_ _00435_ _00408_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12013__A2 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5029_ MuI._0771_ MuI._0772_ MuI._0774_ vssd1 vssd1 vccd1 vccd1 MuI._0775_ sky130_fd_sc_hd__nand3_1
XFILLER_146_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ net132 vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__buf_4
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11772__A1 _00289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11772__B2 _00290_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07066_ _04133_ _06067_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and2_1
XFILLER_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08798__D _00267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__B1 _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._1241__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07968_ _00579_ _00584_ _00564_ _00585_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a211oi_1
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06896__A _04305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09272__A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06919_ _04553_ vssd1 vssd1 vccd1 vccd1 MuI.a_operand\[9\] sky130_fd_sc_hd__clkbuf_2
X_09707_ _06503_ _04100_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__and2_1
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10236__B_N _03680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07899_ _00515_ _00516_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__and2b_1
XANTENNA__10849__C _05025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ _02274_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._4544__B MuI._0603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__D _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09569_ _02195_ _02196_ _02200_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__nand3_1
XANTENNA__08939__A1_N _02851_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11600_ _00444_ _05520_ _04387_ _04388_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__a22o_1
XFILLER_169_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _05275_ _05283_ _05282_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__a21o_1
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10263__A1 _02935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _03295_ _03661_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__and3_1
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13241__B _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._155_ FuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 FuI.Integer\[25\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__11042__A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ _04237_ _04238_ _04239_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21o_1
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ _03626_ _05906_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nand2_2
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFuI._086_ FuI._046_ FuI._049_ FuI.a_operand\[5\] vssd1 vssd1 vccd1 vccd1 FuI._017_
+ sky130_fd_sc_hd__o21a_1
X_10413_ _03108_ _03111_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11977__A _03152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0840_ net132 net116 vssd1 vssd1 vccd1 vccd1 AuI._0060_ sky130_fd_sc_hd__and2b_1
XFILLER_164_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11393_ _02496_ _04391_ _02722_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__o21a_1
XANTENNA_MuI._3607__C MuI._1043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12960__B1 _02731_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _06032_ _06033_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
XANTENNA_input62_A b_operand[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _03019_ _03020_ _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o21a_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09708__A1 _02334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09708__B2 _01332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13063_ _05886_ _05955_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10275_ _06444_ _06442_ _00301_ _04305_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__and4_1
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10318__A2 _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _03432_ _06517_ _06518_ _00278_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__a22o_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10105__B _05467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13268__A1 _03755_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1323_ AuI._0437_ AuI._0517_ AuI._0518_ AuI._0519_ vssd1 vssd1 vccd1 vccd1 AuI._0520_
+ sky130_fd_sc_hd__and4_1
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4400_ MuI._0082_ MuI._3352_ vssd1 vssd1 vccd1 vccd1 MuI._0083_ sky130_fd_sc_hd__xnor2_1
XANTENNA_MuI._4735__A MuI._0321_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5380_ MuI._1158_ MuI._1159_ MuI._1160_ vssd1 vssd1 vccd1 vccd1 MuI._1161_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12916_ _03615_ _05585_ _05660_ _03550_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__a22oi_1
XFILLER_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1254_ AuI._0437_ AuI._0452_ AuI._0453_ AuI._0454_ vssd1 vssd1 vccd1 vccd1 AuI._0456_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10121__A _02916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07498__A2 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4331_ MuI._3294_ MuI._0007_ vssd1 vssd1 vccd1 vccd1 MuI._0008_ sky130_fd_sc_hd__or2_1
XANTENNA_AuI.pe._822__A AuI.operand_a\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _05728_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__xnor2_1
XAuI._1185_ AuI._0389_ AuI._0276_ AuI._0390_ AuI._0212_ vssd1 vssd1 vccd1 vccd1 AuI._0391_
+ sky130_fd_sc_hd__a31o_1
XANTENNA_MuI._5269__C MuI._0017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._4262_ MuI.a_operand\[6\] vssd1 vssd1 vccd1 vccd1 MuI._3362_ sky130_fd_sc_hd__clkbuf_4
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13440__A1 _03842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6001_ MuI._3110_ MuI._3109_ vssd1 vssd1 vccd1 vccd1 MuI._1844_ sky130_fd_sc_hd__and2b_1
XFILLER_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12778_ _05653_ _05654_ _05553_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a21oi_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08526__A _03217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07430__A _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4193_ MuI._3282_ MuI._3284_ vssd1 vssd1 vccd1 vccd1 MuI._3293_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11729_ _00124_ _00125_ _05252_ _05316_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__and4_1
XANTENNA__10494__C _04714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__B1 _00421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12951__B1 _03133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09357__A _02096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08261__A _00877_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._0969_ net118 net14 AuI._0178_ vssd1 vssd1 vccd1 vccd1 AuI._0181_ sky130_fd_sc_hd__mux2_1
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6834_ MuI._2749_ vssd1 vssd1 vccd1 vccd1 MuI.result\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_143_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ _01248_ _01557_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__nor2_1
XFILLER_124_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6765_ MuI._2577_ MuI._2580_ MuI._2587_ vssd1 vssd1 vccd1 vccd1 MuI._2685_ sky130_fd_sc_hd__nand3_2
XFILLER_130_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3977_ MuI._2992_ MuI._2993_ MuI._2990_ MuI._2991_ vssd1 vssd1 vccd1 vccd1 MuI._3077_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08871_ _06503_ _06504_ _06580_ _06581_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__and4_1
XANTENNA__07308__C _06608_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07186__A1 _06470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5716_ MuI._1528_ MuI._1529_ MuI._1526_ vssd1 vssd1 vccd1 vccd1 MuI._1531_ sky130_fd_sc_hd__o21ai_1
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07822_ _00228_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6696_ MuI._2004_ MuI._0793_ MuI._1841_ vssd1 vssd1 vccd1 vccd1 MuI._2609_ sky130_fd_sc_hd__and3b_1
XFILLER_111_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5647_ MuI._1287_ MuI._1331_ vssd1 vssd1 vccd1 vccd1 MuI._1455_ sky130_fd_sc_hd__nand2_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07753_ _00252_ _00212_ _00213_ _00251_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__nand4_1
XAuI.pe._527_ AuI.pe._399_ vssd1 vssd1 vccd1 vccd1 AuI.pe._086_ sky130_fd_sc_hd__buf_2
X_06704_ net111 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__buf_4
XMuI._5578_ MuI._2886_ MuI._0245_ vssd1 vssd1 vccd1 vccd1 MuI._1379_ sky130_fd_sc_hd__nand2_1
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07684_ _03282_ _04176_ _00301_ _00124_ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a22oi_1
XFILLER_71_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XAuI.pe._458_ AuI.pe._022_ vssd1 vssd1 vccd1 vccd1 AuI.pe._023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4529_ MuI._0092_ MuI._0224_ vssd1 vssd1 vccd1 vccd1 MuI._0225_ sky130_fd_sc_hd__nand2_1
X_09423_ _06504_ _00072_ _04434_ _06503_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a22oi_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08139__C _05370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__A1 _00727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__B2 _00728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10966__A net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09354_ _01933_ _01932_ _01931_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__o21ai_1
XFILLER_197_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13431__A1 _05853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _00133_ _00132_ _04240_ _04305_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__and4_1
XANTENNA__13061__B _05660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09285_ _06593_ _00272_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__nand2_1
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08155__B _00398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08236_ _06622_ _04832_ _04896_ _00414_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__a22oi_2
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13195__B1 _03507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ net128 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__buf_2
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07949__B1 _00566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _05788_ _06414_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and2_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _00217_ _00216_ _06591_ _05036_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__nand4_1
XANTENNA__08171__A net29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07049_ _05948_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__buf_4
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6100__A MuI._2791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09714__B _04165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07515__A net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09433__C _00271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__B _06491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _03658_ _04456_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__nand2_1
X_12701_ _02607_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nand2_1
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10893_ _03445_ _03625_ _03627_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand3_1
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _05493_ _05494_ _05495_ _05497_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__o211a_1
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _00676_ _03047_ _06477_ _06444_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__a22oi_1
XFILLER_184_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _04250_ _04252_ _04293_ _04295_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a22oi_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _04872_ _04998_ _05350_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__and4bb_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFuI._138_ FuI._000_ net144 vssd1 vssd1 vccd1 vccd1 FuI.Integer\[9\] sky130_fd_sc_hd__dlxtn_1
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _04067_ _04187_ _04220_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__a211o_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._069_ FuI.a_operand\[25\] vssd1 vssd1 vccd1 vccd1 FuI._037_ sky130_fd_sc_hd__clkbuf_2
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XAuI._0823_ AuI._0040_ AuI._0041_ AuI._0042_ vssd1 vssd1 vccd1 vccd1 AuI._0043_ sky130_fd_sc_hd__and3b_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__xnor2_4
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3900_ MuI.b_operand\[16\] vssd1 vssd1 vccd1 vccd1 MuI._3000_ sky130_fd_sc_hd__clkbuf_2
XFILLER_140_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3634__A MuI._2319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4880_ MuI._0589_ MuI._0590_ MuI._0609_ MuI._0610_ vssd1 vssd1 vccd1 vccd1 MuI._0611_
+ sky130_fd_sc_hd__or4bb_1
X_10327_ _03016_ _03017_ _03018_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__and3_1
X_13115_ _03626_ _05777_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__and2_2
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._6010__A MuI._2550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3831_ MuI._1802_ MuI._2671_ MuI._2440_ MuI._1307_ vssd1 vssd1 vccd1 vccd1 MuI._2931_
+ sky130_fd_sc_hd__a22o_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _03400_ _05970_ _05869_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and3_1
X_10258_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6550_ MuI._2437_ MuI._2447_ vssd1 vssd1 vccd1 vccd1 MuI._2448_ sky130_fd_sc_hd__nor2_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3762_ MuI._2726_ MuI._2715_ vssd1 vssd1 vccd1 vccd1 MuI._2862_ sky130_fd_sc_hd__and2b_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10189_ _02723_ _04671_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__and2b_1
XMuI._5501_ MuI._1292_ MuI._1293_ vssd1 vssd1 vccd1 vccd1 MuI._1294_ sky130_fd_sc_hd__nor2_1
XANTENNA_MuI._5827__A1 MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._6481_ MuI._2368_ MuI._2370_ vssd1 vssd1 vccd1 vccd1 MuI._2372_ sky130_fd_sc_hd__xnor2_1
XMuI._3693_ MuI._2788_ MuI._2792_ vssd1 vssd1 vccd1 vccd1 MuI._2793_ sky130_fd_sc_hd__nor2_1
XMuI._5432_ MuI._1203_ MuI._1205_ vssd1 vssd1 vccd1 vccd1 MuI._1218_ sky130_fd_sc_hd__or2b_1
XAuI._1306_ AuI._0498_ AuI._0499_ AuI._0500_ vssd1 vssd1 vccd1 vccd1 AuI._0504_ sky130_fd_sc_hd__nor3_1
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MuI._3800__C MuI._2867_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5363_ MuI._1077_ MuI._1075_ vssd1 vssd1 vccd1 vccd1 MuI._1143_ sky130_fd_sc_hd__and2b_1
XFILLER_207_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1237_ AuI._0422_ AuI._0439_ vssd1 vssd1 vccd1 vccd1 AuI._0440_ sky130_fd_sc_hd__nand2_1
XANTENNA__11672__B1 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4314_ MuI._3274_ MuI._3273_ vssd1 vssd1 vccd1 vccd1 MuI._3414_ sky130_fd_sc_hd__or2b_1
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5294_ MuI._1063_ MuI._1066_ vssd1 vssd1 vccd1 vccd1 MuI._1067_ sky130_fd_sc_hd__and2_1
XFILLER_179_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1168_ AuI._0262_ AuI._0330_ AuI._0374_ vssd1 vssd1 vccd1 vccd1 AuI._0375_ sky130_fd_sc_hd__or3_4
XFILLER_188_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._4245_ MuI._3342_ MuI._3343_ MuI._3344_ vssd1 vssd1 vccd1 vccd1 MuI._3345_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07160__A net22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._5296__A MuI._0085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XAuI._1099_ AuI._0153_ AuI._0306_ AuI._0308_ AuI._0212_ vssd1 vssd1 vccd1 vccd1 AuI._0309_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11975__A1 _00462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4176_ MuI._3165_ MuI._3258_ MuI._3275_ vssd1 vssd1 vccd1 vccd1 MuI._3276_ sky130_fd_sc_hd__a21o_1
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09070_ _06488_ _06611_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__nand2_1
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11975__B2 _00237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__A1 _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__B2 _02107_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _06511_ _06512_ _06532_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__a21oi_2
XFILLER_129_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3544__A MuI._1285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _02635_ _02636_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__nand2_1
XFILLER_104_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._6817_ MuI._2739_ vssd1 vssd1 vccd1 vccd1 MuI.result\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08923_ _06560_ _04789_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nand2_1
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__B1 _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._6748_ MuI._2656_ MuI._2661_ MuI._2665_ vssd1 vssd1 vccd1 vccd1 MuI._2666_ sky130_fd_sc_hd__and3_1
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08854_ _02539_ _04596_ _01339_ _01338_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a31o_1
XFILLER_57_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12241__A _06444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11565__A2_N _02728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMuI._6679_ MuI._0147_ MuI._2589_ vssd1 vssd1 vccd1 vccd1 MuI._2590_ sky130_fd_sc_hd__xnor2_1
X_07805_ _05112_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__buf_4
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _01388_ _01393_ _01402_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__a21oi_4
XFILLER_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07736_ _00129_ _00139_ _00138_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a21o_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_AuI.pe._462__A AuI.pe._024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ _00280_ _00284_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__nor2_2
XANTENNA_MuI._6243__A1 MuI._1153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._6243__B2 MuI._0735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__B2 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__A _03809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09406_ _02012_ _02014_ _02023_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__and3_1
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07598_ _00029_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__buf_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07070__A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09337_ _01952_ _01953_ _01954_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__nand3_1
XANTENNA__11304__B _03282_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4006__B1 MuI._2797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ net108 _00098_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__nand2_1
XANTENNA__10086__A_N _02388_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08219_ _02528_ _05036_ _00537_ _00538_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _06460_ _04703_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__nand2_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11718__A1 _00058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ _03904_ _03905_ _03989_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__nand4_4
XFILLER_181_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_MuI._3454__A MuI._0339_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11161_ _03912_ _03915_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__and2_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07229__B _06529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__A2 _06056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _04542_ _02604_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__or2b_1
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ _04262_ _02728_ _03675_ _04327_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ _02118_ _03917_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__or2b_1
XFILLER_209_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07890__D _00287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_AuI._0946__A0 net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07245__A _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A a_operand[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4493__B1 MuI._2845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__B1 _03971_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ _04810_ _04812_ _04700_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _02345_ _04197_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__or2b_1
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1022_ AuI._0223_ AuI._0225_ AuI._0227_ AuI._0231_ AuI._0233_ vssd1 vssd1 vccd1
+ vccd1 AuI._0234_ sky130_fd_sc_hd__o311a_1
XFILLER_204_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI._0855__A_N net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _03606_ _03607_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__or3_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11214__B _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _05480_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and2b_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._4030_ MuI._0570_ MuI._2975_ MuI._2976_ MuI._0339_ vssd1 vssd1 vccd1 vccd1 MuI._3130_
+ sky130_fd_sc_hd__a22o_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12546_ _00133_ _00132_ _05884_ _00789_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__nand4_1
XANTENNA__08822__A1 _00150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08822__B2 _06494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12477_ _05289_ _05290_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and4_1
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08523__B _01140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5981_ MuI._1819_ MuI._1821_ vssd1 vssd1 vccd1 vccd1 MuI._1822_ sky130_fd_sc_hd__xor2_2
XANTENNA_output93_A net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11428_ _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__nor2_1
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11587__D _00783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4932_ MuI._0664_ MuI._0665_ vssd1 vssd1 vccd1 vccd1 MuI._0668_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._0806_ net18 vssd1 vssd1 vccd1 vccd1 AuI._0026_ sky130_fd_sc_hd__inv_2
X_11359_ _04127_ _04128_ _03888_ _03892_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o211ai_1
XFILLER_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI.pe._792_ AuI.pe._393_ AuI.pe._105_ AuI.pe._380_ AuI.pe._149_ AuI.pe._395_ vssd1
+ vssd1 vccd1 vccd1 AuI.pe._332_ sky130_fd_sc_hd__o311a_1
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._4863_ MuI._2838_ MuI._2765_ MuI._2785_ MuI._2836_ vssd1 vssd1 vccd1 vccd1 MuI._0593_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6602_ MuI._0999_ MuI._2482_ MuI._2483_ vssd1 vssd1 vccd1 vccd1 MuI._2505_ sky130_fd_sc_hd__nor3_4
XFILLER_141_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._3814_ MuI._2682_ vssd1 vssd1 vccd1 vccd1 MuI._2914_ sky130_fd_sc_hd__buf_2
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4794_ MuI._0510_ MuI._0514_ MuI._0516_ vssd1 vssd1 vccd1 vccd1 MuI._0517_ sky130_fd_sc_hd__o21ai_2
X_13029_ _02639_ _05843_ _01847_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__o21ai_4
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08896__D _00030_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6533_ MuI._2228_ MuI._2428_ vssd1 vssd1 vccd1 vccd1 MuI._2430_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMuI._3745_ MuI._2837_ vssd1 vssd1 vccd1 vccd1 MuI._2845_ sky130_fd_sc_hd__clkbuf_4
XFILLER_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07155__A _03561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._6464_ MuI._1962_ MuI._1980_ vssd1 vssd1 vccd1 vccd1 MuI._2354_ sky130_fd_sc_hd__or2b_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._3676_ MuI.a_operand\[10\] vssd1 vssd1 vccd1 vccd1 MuI._2765_ sky130_fd_sc_hd__buf_2
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _01135_ _01174_ _01186_ _01187_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__o211a_2
XANTENNA_MuI._4484__B1 MuI._0175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06994__A net19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._5415_ MuI._1192_ MuI._1193_ MuI._1198_ vssd1 vssd1 vccd1 vccd1 MuI._1200_ sky130_fd_sc_hd__nand3_1
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09370__A _02420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _00135_ _00136_ _00137_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a21o_1
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._6395_ MuI._2251_ MuI._2267_ MuI._2274_ MuI._2277_ vssd1 vssd1 vccd1 vccd1 MuI._2278_
+ sky130_fd_sc_hd__a211o_1
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._5346_ MuI._2892_ MuI._2319_ MuI._3185_ MuI._2829_ vssd1 vssd1 vccd1 vccd1 MuI._1124_
+ sky130_fd_sc_hd__and4_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ _00044_ _00055_ _00068_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07602__B _06613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13398__B1 _02745_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3539__A MuI._1274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5277_ MuI._1030_ MuI._1046_ MuI._1047_ vssd1 vssd1 vccd1 vccd1 MuI._1048_ sky130_fd_sc_hd__nand3_2
XANTENNA__10666__D _06568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ _06682_ _06525_ _06568_ _00000_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_188_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4228_ MuI._2616_ MuI._2660_ MuI._2844_ MuI._2845_ vssd1 vssd1 vccd1 vccd1 MuI._3328_
+ sky130_fd_sc_hd__and4_1
X_09122_ _02851_ _04057_ _01738_ _01739_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a31o_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08714__A net110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMuI._4159_ MuI._3195_ MuI._3188_ MuI._3194_ vssd1 vssd1 vccd1 vccd1 MuI._3259_ sky130_fd_sc_hd__and3_1
XFILLER_136_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09053_ _01669_ _01670_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nor2_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07975__D _00089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _06508_ _06498_ _06507_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__nand3_1
XFILLER_190_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09369__A2 _00592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10384__B1 _00153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09955_ _02617_ _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__xor2_2
XANTENNA_MuI._6585__A MuI._2486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._4850__A1_N MuI._2451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _01522_ _01523_ _06608_ _00259_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__and4bb_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _02538_ _02542_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__o21a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_AuI._0928__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _01444_ _01442_ _01443_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__or3_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _01384_ _01385_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__and2b_1
XANTENNA__07917__A1_N _02528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10439__A1 _02977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07719_ _06455_ _06456_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__nor2_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08699_ _01275_ _01315_ _01316_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__a21bo_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._4227__B1 MuI._2976_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ _02229_ _00385_ _05820_ _02431_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a22o_1
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07512__B _00081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _03337_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__xor2_1
XFILLER_186_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _04929_ _02727_ _05249_ _04011_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12061__B1 _04642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ _06237_ _06241_ _06291_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__nor3_1
X_10592_ _02767_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__o21a_1
XFILLER_194_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _05158_ _05173_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and2_1
XANTENNA__12146__A _04956_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12262_ _04962_ _04964_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nand2_1
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09158__C _00082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__A1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFuI._142__148 vssd1 vssd1 vccd1 vccd1 FuI._142__148/HI net148 sky130_fd_sc_hd__conb_1
XFILLER_123_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _00081_ _05187_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__and2_2
XFILLER_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XAuI._1640_ AuI._0802_ AuI._0803_ vssd1 vssd1 vccd1 vccd1 AuI._0804_ sky130_fd_sc_hd__and2_1
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12193_ MuI.result\[14\] _02739_ _03494_ _02795_ _05026_ vssd1 vssd1 vccd1 vccd1
+ _05027_ sky130_fd_sc_hd__a221o_1
XFILLER_150_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11144_ _03727_ _03880_ _03896_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__o211ai_2
XAuI._1571_ AuI.pe.Significand\[9\] AuI._0721_ vssd1 vssd1 vccd1 vccd1 AuI._0748_
+ sky130_fd_sc_hd__or2_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 ALU_Output[14] sky130_fd_sc_hd__buf_2
XFILLER_110_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 ALU_Output[24] sky130_fd_sc_hd__buf_2
XANTENNA__12116__A1 _00534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 ALU_Output[5] sky130_fd_sc_hd__buf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MuI._3912__A MuI._2817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _03696_ _03823_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__xor2_4
XFILLER_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ _01328_ _01329_ _00954_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11209__B _03099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._3530_ MuI._1164_ MuI._0526_ MuI._0757_ vssd1 vssd1 vccd1 vccd1 MuI._1186_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12419__A2 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMuI._3461_ MuI._0405_ MuI._0416_ vssd1 vssd1 vccd1 vccd1 MuI._0427_ sky130_fd_sc_hd__or2_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__A _00292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5200_ MuI._0798_ MuI._0962_ vssd1 vssd1 vccd1 vccd1 MuI._0963_ sky130_fd_sc_hd__nor2_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11977_ _03152_ _00398_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__nand2_1
XMuI._6180_ MuI._2034_ MuI._2039_ MuI._2040_ vssd1 vssd1 vccd1 vccd1 MuI._2041_ sky130_fd_sc_hd__nand3_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10928_ _02703_ _03295_ _03661_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a31oi_1
XFILLER_177_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._5131_ MuI._2871_ MuI._0101_ vssd1 vssd1 vccd1 vccd1 MuI._0887_ sky130_fd_sc_hd__nand2_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_AuI.pe._830__A AuI.operand_a\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XAuI._1005_ AuI._0190_ AuI._0191_ AuI._0216_ vssd1 vssd1 vccd1 vccd1 AuI._0217_ sky130_fd_sc_hd__or3b_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ _03588_ _03571_ _03573_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__and3_1
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMuI._5062_ MuI._0807_ MuI._0810_ vssd1 vssd1 vccd1 vccd1 MuI._0811_ sky130_fd_sc_hd__nor2_1
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08534__A _00915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._4013_ MuI._3112_ vssd1 vssd1 vccd1 vccd1 MuI._3113_ sky130_fd_sc_hd__inv_2
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MuI._3992__A2 MuI._2860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _02970_ _04994_ _05375_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09349__B _06480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XMuI._5964_ MuI._1798_ MuI._1801_ MuI._1803_ vssd1 vssd1 vccd1 vccd1 MuI._1804_ sky130_fd_sc_hd__and3_1
XFILLER_126_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A _05305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4915_ MuI._0455_ MuI._0648_ MuI._0609_ MuI._0607_ vssd1 vssd1 vccd1 vccd1 MuI._0650_
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__09365__A _06663_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMuI._5895_ MuI._1727_ vssd1 vssd1 vccd1 vccd1 MuI._1728_ sky130_fd_sc_hd__inv_2
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMuI._4846_ MuI.a_operand\[13\] MuI.a_operand\[12\] MuI._2866_ MuI._2868_ vssd1 vssd1
+ vccd1 vccd1 MuI._0574_ sky130_fd_sc_hd__and4_1
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _02309_ _02311_ _02310_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09084__B _00093_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06952_ _04907_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__clkbuf_8
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

