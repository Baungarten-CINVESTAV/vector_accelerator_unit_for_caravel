magic
tech sky130A
magscale 1 2
timestamp 1669389075
<< obsli1 >>
rect 1104 2159 98808 117521
<< obsm1 >>
rect 14 1300 99898 117552
<< metal2 >>
rect 2594 119200 2650 119800
rect 6458 119200 6514 119800
rect 10322 119200 10378 119800
rect 14830 119200 14886 119800
rect 18694 119200 18750 119800
rect 23202 119200 23258 119800
rect 27066 119200 27122 119800
rect 31574 119200 31630 119800
rect 35438 119200 35494 119800
rect 39946 119200 40002 119800
rect 43810 119200 43866 119800
rect 48318 119200 48374 119800
rect 52182 119200 52238 119800
rect 56690 119200 56746 119800
rect 60554 119200 60610 119800
rect 65062 119200 65118 119800
rect 68926 119200 68982 119800
rect 72790 119200 72846 119800
rect 77298 119200 77354 119800
rect 81162 119200 81218 119800
rect 85670 119200 85726 119800
rect 89534 119200 89590 119800
rect 94042 119200 94098 119800
rect 97906 119200 97962 119800
rect 18 200 74 800
rect 3882 200 3938 800
rect 7746 200 7802 800
rect 12254 200 12310 800
rect 16118 200 16174 800
rect 20626 200 20682 800
rect 24490 200 24546 800
rect 28998 200 29054 800
rect 32862 200 32918 800
rect 37370 200 37426 800
rect 41234 200 41290 800
rect 45742 200 45798 800
rect 49606 200 49662 800
rect 54114 200 54170 800
rect 57978 200 58034 800
rect 61842 200 61898 800
rect 66350 200 66406 800
rect 70214 200 70270 800
rect 74722 200 74778 800
rect 78586 200 78642 800
rect 83094 200 83150 800
rect 86958 200 87014 800
rect 91466 200 91522 800
rect 95330 200 95386 800
rect 99838 200 99894 800
<< obsm2 >>
rect 20 119856 99892 119898
rect 20 119144 2538 119856
rect 2706 119144 6402 119856
rect 6570 119144 10266 119856
rect 10434 119144 14774 119856
rect 14942 119144 18638 119856
rect 18806 119144 23146 119856
rect 23314 119144 27010 119856
rect 27178 119144 31518 119856
rect 31686 119144 35382 119856
rect 35550 119144 39890 119856
rect 40058 119144 43754 119856
rect 43922 119144 48262 119856
rect 48430 119144 52126 119856
rect 52294 119144 56634 119856
rect 56802 119144 60498 119856
rect 60666 119144 65006 119856
rect 65174 119144 68870 119856
rect 69038 119144 72734 119856
rect 72902 119144 77242 119856
rect 77410 119144 81106 119856
rect 81274 119144 85614 119856
rect 85782 119144 89478 119856
rect 89646 119144 93986 119856
rect 94154 119144 97850 119856
rect 98018 119144 99892 119856
rect 20 856 99892 119144
rect 130 800 3826 856
rect 3994 800 7690 856
rect 7858 800 12198 856
rect 12366 800 16062 856
rect 16230 800 20570 856
rect 20738 800 24434 856
rect 24602 800 28942 856
rect 29110 800 32806 856
rect 32974 800 37314 856
rect 37482 800 41178 856
rect 41346 800 45686 856
rect 45854 800 49550 856
rect 49718 800 54058 856
rect 54226 800 57922 856
rect 58090 800 61786 856
rect 61954 800 66294 856
rect 66462 800 70158 856
rect 70326 800 74666 856
rect 74834 800 78530 856
rect 78698 800 83038 856
rect 83206 800 86902 856
rect 87070 800 91410 856
rect 91578 800 95274 856
rect 95442 800 99782 856
<< metal3 >>
rect 200 118328 800 118448
rect 99200 117648 99800 117768
rect 200 114248 800 114368
rect 99200 113568 99800 113688
rect 200 109488 800 109608
rect 99200 108808 99800 108928
rect 200 105408 800 105528
rect 99200 104728 99800 104848
rect 200 100648 800 100768
rect 99200 99968 99800 100088
rect 200 96568 800 96688
rect 99200 95888 99800 96008
rect 200 91808 800 91928
rect 99200 91128 99800 91248
rect 200 87728 800 87848
rect 99200 87048 99800 87168
rect 200 82968 800 83088
rect 99200 82968 99800 83088
rect 200 78888 800 79008
rect 99200 78208 99800 78328
rect 200 74128 800 74248
rect 99200 74128 99800 74248
rect 200 70048 800 70168
rect 99200 69368 99800 69488
rect 200 65288 800 65408
rect 99200 65288 99800 65408
rect 200 61208 800 61328
rect 99200 60528 99800 60648
rect 200 57128 800 57248
rect 99200 56448 99800 56568
rect 200 52368 800 52488
rect 99200 51688 99800 51808
rect 200 48288 800 48408
rect 99200 47608 99800 47728
rect 200 43528 800 43648
rect 99200 42848 99800 42968
rect 200 39448 800 39568
rect 99200 38768 99800 38888
rect 200 34688 800 34808
rect 99200 34008 99800 34128
rect 200 30608 800 30728
rect 99200 29928 99800 30048
rect 200 25848 800 25968
rect 99200 25168 99800 25288
rect 200 21768 800 21888
rect 99200 21088 99800 21208
rect 200 17008 800 17128
rect 99200 17008 99800 17128
rect 200 12928 800 13048
rect 99200 12248 99800 12368
rect 200 8168 800 8288
rect 99200 8168 99800 8288
rect 200 4088 800 4208
rect 99200 3408 99800 3528
<< obsm3 >>
rect 880 118248 99200 118421
rect 565 117848 99200 118248
rect 565 117568 99120 117848
rect 565 114448 99200 117568
rect 880 114168 99200 114448
rect 565 113768 99200 114168
rect 565 113488 99120 113768
rect 565 109688 99200 113488
rect 880 109408 99200 109688
rect 565 109008 99200 109408
rect 565 108728 99120 109008
rect 565 105608 99200 108728
rect 880 105328 99200 105608
rect 565 104928 99200 105328
rect 565 104648 99120 104928
rect 565 100848 99200 104648
rect 880 100568 99200 100848
rect 565 100168 99200 100568
rect 565 99888 99120 100168
rect 565 96768 99200 99888
rect 880 96488 99200 96768
rect 565 96088 99200 96488
rect 565 95808 99120 96088
rect 565 92008 99200 95808
rect 880 91728 99200 92008
rect 565 91328 99200 91728
rect 565 91048 99120 91328
rect 565 87928 99200 91048
rect 880 87648 99200 87928
rect 565 87248 99200 87648
rect 565 86968 99120 87248
rect 565 83168 99200 86968
rect 880 82888 99120 83168
rect 565 79088 99200 82888
rect 880 78808 99200 79088
rect 565 78408 99200 78808
rect 565 78128 99120 78408
rect 565 74328 99200 78128
rect 880 74048 99120 74328
rect 565 70248 99200 74048
rect 880 69968 99200 70248
rect 565 69568 99200 69968
rect 565 69288 99120 69568
rect 565 65488 99200 69288
rect 880 65208 99120 65488
rect 565 61408 99200 65208
rect 880 61128 99200 61408
rect 565 60728 99200 61128
rect 565 60448 99120 60728
rect 565 57328 99200 60448
rect 880 57048 99200 57328
rect 565 56648 99200 57048
rect 565 56368 99120 56648
rect 565 52568 99200 56368
rect 880 52288 99200 52568
rect 565 51888 99200 52288
rect 565 51608 99120 51888
rect 565 48488 99200 51608
rect 880 48208 99200 48488
rect 565 47808 99200 48208
rect 565 47528 99120 47808
rect 565 43728 99200 47528
rect 880 43448 99200 43728
rect 565 43048 99200 43448
rect 565 42768 99120 43048
rect 565 39648 99200 42768
rect 880 39368 99200 39648
rect 565 38968 99200 39368
rect 565 38688 99120 38968
rect 565 34888 99200 38688
rect 880 34608 99200 34888
rect 565 34208 99200 34608
rect 565 33928 99120 34208
rect 565 30808 99200 33928
rect 880 30528 99200 30808
rect 565 30128 99200 30528
rect 565 29848 99120 30128
rect 565 26048 99200 29848
rect 880 25768 99200 26048
rect 565 25368 99200 25768
rect 565 25088 99120 25368
rect 565 21968 99200 25088
rect 880 21688 99200 21968
rect 565 21288 99200 21688
rect 565 21008 99120 21288
rect 565 17208 99200 21008
rect 880 16928 99120 17208
rect 565 13128 99200 16928
rect 880 12848 99200 13128
rect 565 12448 99200 12848
rect 565 12168 99120 12448
rect 565 8368 99200 12168
rect 880 8088 99120 8368
rect 565 4288 99200 8088
rect 880 4008 99200 4288
rect 565 3608 99200 4008
rect 565 3328 99120 3608
rect 565 1939 99200 3328
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
<< obsm4 >>
rect 979 2048 4128 117197
rect 4608 2048 19488 117197
rect 19968 2048 34848 117197
rect 35328 2048 50208 117197
rect 50688 2048 65568 117197
rect 66048 2048 80928 117197
rect 81408 2048 89181 117197
rect 979 1939 89181 2048
<< labels >>
rlabel metal3 s 200 57128 800 57248 6 ALU_Output[0]
port 1 nsew signal output
rlabel metal2 s 28998 200 29054 800 6 ALU_Output[10]
port 2 nsew signal output
rlabel metal3 s 99200 91128 99800 91248 6 ALU_Output[11]
port 3 nsew signal output
rlabel metal3 s 99200 29928 99800 30048 6 ALU_Output[12]
port 4 nsew signal output
rlabel metal3 s 99200 117648 99800 117768 6 ALU_Output[13]
port 5 nsew signal output
rlabel metal3 s 99200 42848 99800 42968 6 ALU_Output[14]
port 6 nsew signal output
rlabel metal3 s 200 105408 800 105528 6 ALU_Output[15]
port 7 nsew signal output
rlabel metal3 s 200 100648 800 100768 6 ALU_Output[16]
port 8 nsew signal output
rlabel metal2 s 60554 119200 60610 119800 6 ALU_Output[17]
port 9 nsew signal output
rlabel metal2 s 94042 119200 94098 119800 6 ALU_Output[18]
port 10 nsew signal output
rlabel metal3 s 200 48288 800 48408 6 ALU_Output[19]
port 11 nsew signal output
rlabel metal3 s 99200 25168 99800 25288 6 ALU_Output[1]
port 12 nsew signal output
rlabel metal3 s 200 82968 800 83088 6 ALU_Output[20]
port 13 nsew signal output
rlabel metal2 s 91466 200 91522 800 6 ALU_Output[21]
port 14 nsew signal output
rlabel metal3 s 200 12928 800 13048 6 ALU_Output[22]
port 15 nsew signal output
rlabel metal3 s 99200 104728 99800 104848 6 ALU_Output[23]
port 16 nsew signal output
rlabel metal2 s 61842 200 61898 800 6 ALU_Output[24]
port 17 nsew signal output
rlabel metal2 s 12254 200 12310 800 6 ALU_Output[25]
port 18 nsew signal output
rlabel metal3 s 200 70048 800 70168 6 ALU_Output[26]
port 19 nsew signal output
rlabel metal2 s 95330 200 95386 800 6 ALU_Output[27]
port 20 nsew signal output
rlabel metal3 s 99200 113568 99800 113688 6 ALU_Output[28]
port 21 nsew signal output
rlabel metal2 s 85670 119200 85726 119800 6 ALU_Output[29]
port 22 nsew signal output
rlabel metal3 s 200 74128 800 74248 6 ALU_Output[2]
port 23 nsew signal output
rlabel metal3 s 200 25848 800 25968 6 ALU_Output[30]
port 24 nsew signal output
rlabel metal2 s 45742 200 45798 800 6 ALU_Output[31]
port 25 nsew signal output
rlabel metal3 s 99200 95888 99800 96008 6 ALU_Output[3]
port 26 nsew signal output
rlabel metal3 s 99200 65288 99800 65408 6 ALU_Output[4]
port 27 nsew signal output
rlabel metal3 s 99200 69368 99800 69488 6 ALU_Output[5]
port 28 nsew signal output
rlabel metal2 s 56690 119200 56746 119800 6 ALU_Output[6]
port 29 nsew signal output
rlabel metal3 s 99200 82968 99800 83088 6 ALU_Output[7]
port 30 nsew signal output
rlabel metal3 s 200 52368 800 52488 6 ALU_Output[8]
port 31 nsew signal output
rlabel metal3 s 200 78888 800 79008 6 ALU_Output[9]
port 32 nsew signal output
rlabel metal2 s 27066 119200 27122 119800 6 Exception
port 33 nsew signal output
rlabel metal3 s 99200 108808 99800 108928 6 Operation[0]
port 34 nsew signal input
rlabel metal2 s 31574 119200 31630 119800 6 Operation[1]
port 35 nsew signal input
rlabel metal2 s 52182 119200 52238 119800 6 Operation[2]
port 36 nsew signal input
rlabel metal3 s 99200 47608 99800 47728 6 Operation[3]
port 37 nsew signal input
rlabel metal2 s 35438 119200 35494 119800 6 Overflow
port 38 nsew signal output
rlabel metal2 s 18694 119200 18750 119800 6 Underflow
port 39 nsew signal output
rlabel metal2 s 48318 119200 48374 119800 6 a_operand[0]
port 40 nsew signal input
rlabel metal2 s 24490 200 24546 800 6 a_operand[10]
port 41 nsew signal input
rlabel metal2 s 39946 119200 40002 119800 6 a_operand[11]
port 42 nsew signal input
rlabel metal3 s 99200 8168 99800 8288 6 a_operand[12]
port 43 nsew signal input
rlabel metal3 s 99200 56448 99800 56568 6 a_operand[13]
port 44 nsew signal input
rlabel metal2 s 68926 119200 68982 119800 6 a_operand[14]
port 45 nsew signal input
rlabel metal2 s 23202 119200 23258 119800 6 a_operand[15]
port 46 nsew signal input
rlabel metal3 s 99200 12248 99800 12368 6 a_operand[16]
port 47 nsew signal input
rlabel metal3 s 99200 99968 99800 100088 6 a_operand[17]
port 48 nsew signal input
rlabel metal3 s 200 87728 800 87848 6 a_operand[18]
port 49 nsew signal input
rlabel metal2 s 78586 200 78642 800 6 a_operand[19]
port 50 nsew signal input
rlabel metal2 s 41234 200 41290 800 6 a_operand[1]
port 51 nsew signal input
rlabel metal3 s 99200 34008 99800 34128 6 a_operand[20]
port 52 nsew signal input
rlabel metal3 s 200 61208 800 61328 6 a_operand[21]
port 53 nsew signal input
rlabel metal3 s 200 8168 800 8288 6 a_operand[22]
port 54 nsew signal input
rlabel metal3 s 99200 3408 99800 3528 6 a_operand[23]
port 55 nsew signal input
rlabel metal3 s 200 21768 800 21888 6 a_operand[24]
port 56 nsew signal input
rlabel metal2 s 83094 200 83150 800 6 a_operand[25]
port 57 nsew signal input
rlabel metal2 s 81162 119200 81218 119800 6 a_operand[26]
port 58 nsew signal input
rlabel metal2 s 70214 200 70270 800 6 a_operand[27]
port 59 nsew signal input
rlabel metal2 s 7746 200 7802 800 6 a_operand[28]
port 60 nsew signal input
rlabel metal2 s 32862 200 32918 800 6 a_operand[29]
port 61 nsew signal input
rlabel metal2 s 99838 200 99894 800 6 a_operand[2]
port 62 nsew signal input
rlabel metal3 s 200 4088 800 4208 6 a_operand[30]
port 63 nsew signal input
rlabel metal3 s 99200 38768 99800 38888 6 a_operand[31]
port 64 nsew signal input
rlabel metal3 s 200 17008 800 17128 6 a_operand[3]
port 65 nsew signal input
rlabel metal3 s 200 91808 800 91928 6 a_operand[4]
port 66 nsew signal input
rlabel metal3 s 99200 17008 99800 17128 6 a_operand[5]
port 67 nsew signal input
rlabel metal2 s 2594 119200 2650 119800 6 a_operand[6]
port 68 nsew signal input
rlabel metal3 s 99200 51688 99800 51808 6 a_operand[7]
port 69 nsew signal input
rlabel metal3 s 99200 78208 99800 78328 6 a_operand[8]
port 70 nsew signal input
rlabel metal2 s 86958 200 87014 800 6 a_operand[9]
port 71 nsew signal input
rlabel metal3 s 99200 87048 99800 87168 6 b_operand[0]
port 72 nsew signal input
rlabel metal2 s 6458 119200 6514 119800 6 b_operand[10]
port 73 nsew signal input
rlabel metal3 s 200 65288 800 65408 6 b_operand[11]
port 74 nsew signal input
rlabel metal2 s 54114 200 54170 800 6 b_operand[12]
port 75 nsew signal input
rlabel metal2 s 18 200 74 800 6 b_operand[13]
port 76 nsew signal input
rlabel metal2 s 66350 200 66406 800 6 b_operand[14]
port 77 nsew signal input
rlabel metal2 s 10322 119200 10378 119800 6 b_operand[15]
port 78 nsew signal input
rlabel metal2 s 43810 119200 43866 119800 6 b_operand[16]
port 79 nsew signal input
rlabel metal3 s 200 34688 800 34808 6 b_operand[17]
port 80 nsew signal input
rlabel metal3 s 200 109488 800 109608 6 b_operand[18]
port 81 nsew signal input
rlabel metal2 s 16118 200 16174 800 6 b_operand[19]
port 82 nsew signal input
rlabel metal2 s 3882 200 3938 800 6 b_operand[1]
port 83 nsew signal input
rlabel metal2 s 89534 119200 89590 119800 6 b_operand[20]
port 84 nsew signal input
rlabel metal2 s 65062 119200 65118 119800 6 b_operand[21]
port 85 nsew signal input
rlabel metal2 s 49606 200 49662 800 6 b_operand[22]
port 86 nsew signal input
rlabel metal2 s 97906 119200 97962 119800 6 b_operand[23]
port 87 nsew signal input
rlabel metal3 s 99200 21088 99800 21208 6 b_operand[24]
port 88 nsew signal input
rlabel metal3 s 200 114248 800 114368 6 b_operand[25]
port 89 nsew signal input
rlabel metal3 s 200 43528 800 43648 6 b_operand[26]
port 90 nsew signal input
rlabel metal2 s 20626 200 20682 800 6 b_operand[27]
port 91 nsew signal input
rlabel metal2 s 37370 200 37426 800 6 b_operand[28]
port 92 nsew signal input
rlabel metal3 s 200 39448 800 39568 6 b_operand[29]
port 93 nsew signal input
rlabel metal3 s 99200 74128 99800 74248 6 b_operand[2]
port 94 nsew signal input
rlabel metal2 s 57978 200 58034 800 6 b_operand[30]
port 95 nsew signal input
rlabel metal2 s 77298 119200 77354 119800 6 b_operand[31]
port 96 nsew signal input
rlabel metal2 s 72790 119200 72846 119800 6 b_operand[3]
port 97 nsew signal input
rlabel metal3 s 200 118328 800 118448 6 b_operand[4]
port 98 nsew signal input
rlabel metal2 s 14830 119200 14886 119800 6 b_operand[5]
port 99 nsew signal input
rlabel metal2 s 74722 200 74778 800 6 b_operand[6]
port 100 nsew signal input
rlabel metal3 s 200 30608 800 30728 6 b_operand[7]
port 101 nsew signal input
rlabel metal3 s 200 96568 800 96688 6 b_operand[8]
port 102 nsew signal input
rlabel metal3 s 99200 60528 99800 60648 6 b_operand[9]
port 103 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 104 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 105 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 45828474
string GDS_FILE /home/baungarten/Caravel_4_ALU/openlane/ALU/runs/22_11_25_09_01/results/signoff/ALU.magic.gds
string GDS_START 1253760
<< end >>

